��   v	�A��*SYST�EM*��V8.3�0340 11�/9/2020 A   ����UI_CON�FIG_T  �� B$NUM�_MENUS � 9* NECT�CRECOVER�>CCOLOR_�CRR:EXTS�TAT��$TO�P>_IDXCMEM_LIMIR�$DBGLVL��POPUP_M�ASK�zA � $DUMMY�63�ODE�
4�CFOCA �5VCPS)C��g �HAN� � T�IMEOU�PI�PESIZE ޡ MWIN�PA�NEMAP�  �� � FAVB ?�� 
$HL�_�DIQ?� qEgLEMZ�UR� �l� Ss�$H�MI�RO+\~W ADONLY� }�TOUCH��PROOMMO�#?$�ALAR�< �FILVEW�	ENB=%%�fC 1"USER�:)FCTN:)WI��� I* _ED��l"V!_TITL�� 1"COOR{DF<#LOCK6%��$F%�!b"EBF�OR�? �"e&
�"�%�!BA�!j ?��"BG�%�!jI{NSR$IO}�7PM�X_PK}T�"IHELP� �MER�BLNK�C=ENAB�!? SIPMANUA�pL4"="�BEEY�?$�=&q!EDy#�M0IP0q!�JWD8�D7�DSB�� �GTB9I�:J�<BT_DEVICg1� &USTOM~0 t $} RT_SPID�r8DC@D*PAG� �?^C\ISCR�EuEF��UGN~�@$FLAG��@�&�1  �h 	$PWD_ACCES� E ��8��C�!�%)�$LABE� $Tz j�@�3
R��	 #BUSRV�I 1  < �`�B*�B� QPR�I�m� t1^PT�RIP�"m�$$�CLA�@ �S��Q��R��RtP�\ SI�}W�  ���QI�RTs1}_�P'2 L�3hL3!x�R	 /,��?����R�P�S�S�Q|�� , �!@yo��
 ���Q�]ooo�o�o�o�o�o  Yo�o $6H�o l~����U� �� �2�D�V��z� ������ԏc���
� �.�@�R��v����� ����П�q���*� <�N�`�������� ̯ޯm���&�8�J��\�n��PTP�TX������{�� s �{���$�/softpar�t/genlin�k?help=/�md/tpmenu.dgp�
��.��@���&տ�pwd ���ϟϱ��������� ��/�A���e�w߉� �߭߿�N�`�����+�=�O�����Qb3ff�St�($�߀���������������Q�Q�o|���� ���Rcz�4a��6�e����  ��L"P����L���z����5��/`  1�b�����  �S)B� 1�XR �\�}!@wREG VED���0wholemod.htmD	�singlUd�oubltr�ip�brows�L�1��� �-?Qc��?Qdev.s�Zl��1�	t/����W/i/ {/E/�/�/�/�/�/?� �P(?:?L?^?�p?�?�?�?�?�?�6 @$?�?O�?/OAOSO "F	??�O�O�O�O �O�O�O__)_;_M_ __q_�_�_�_�_�_� �_�_oo/oAoSoeo wo�o�o�o�o�o�o�o +=O?�� �������,� 'OP�b�1�C�����aO sOY�����:�5� G�Y���}�����ʟş ן�����_?�9� g�y���������ӯ� ��	��-�?�Q�c�u� ������y���
�� .�@�R�d�vψσ��� �ύϟ���߽�Ϗ�� N�I�[�mߖߑߣߵ� ��������&�!�3�E� n�i�{�I�������� ������/�A�S�e� w��������������� տBTfx�� ������� �Pb�+��� �����/:/5/ G/Y/�/}/�/�/�/�/ �/���/�/?1?C?U? g?y?�?�?�?�?�?�? �?	OO-O?OQOcO1 �O�O�O�O�O�O
__ ._@_;d_v_E_W_�_��_�Z�$UI_T�OPMENU 1��P�QR� 
d�QvA)�*defaul�t�OjM*le�vel0 *lK	G  o0coo�aosbtpio[2�3]8tpst[1�huo�o�oCoUo� =
h58E01�.gif8	m�enu56y-pXq1!36zWr5zUt4]{Dq������� �*�uB�S�e�w��������<�prim�=Xqpage,1422,1����� �#�5�@�Y�k�}���衟��B�Ȇclass,5�����h'�9�D�М13@�@v���������E�Ȍ53ڏ����0�B�
E�Ȍ8�}����� ��ſD������1�C�nI�P�Qo{�*m�m�qkϥ�ϭftyx�m�o�amf[0�o���	��c[164�g>�59�hq���{�Qx2�[}��qz} gw5{�߹s[�m�F�X� j�|��ٿ�������� �����0�B�T�f�x����ϝ2�������� ��ڟOas� �&8d���� ϯ�14�^p���%�ȃainedis���//�%/ �confi�g=single}&ȂwintpԀ 0/p/�/�/�/mJ�Qf� �/�/+e�/�o��?/? A?T?e?w?�?�?	?�? �?�?�?OO+O=OOO �qO�O�O�O�O�O�O %�_(_:_L_^_p_�O �_�_�_�_�_�_}_ o $o6oHoZolo~oo�o �o�o�o�o�o�o 2 DVhz	��� ���
��.�@�R� d�v��������Џ���]Nc�<��ϙ� ����iO���s�ͤ�ɟ�ϱ�u��|�f�؟ >�4����Z����ߤ�6��u7���0�	� �-�?�Q���u����� ����Ͽ^����)�P;�M�_�>"41C �ϫϽ�������� )�;�M�_��σߕߧ� ��������2��%�7� I�[�m����6t�����������<$�74 ��-�?�Q�c�u��,�����%	TPTX[�209�,���24`�����Σ��18���������0`2����1o�A�i�tv ������0�
��1�
ӯ�C:D$tr?eeviewQ#��3�&dual=�oe81,26,4����~��� //+/=/�a/s/�/��/�/�/��;P�53p��'?9?K?V/ o?�?�?�?�?�?X?�? �?O#O5OGO�/�/�	1�/�2f��O�O�O� �6hO�edit���O�O,_>_P_�� O�	_S\_�_�_�_ ���_oW�o�-o� Soeowo�o�o�o�o�o ?o�o+=Oa t�㥝���� ���?B�T�f�x��� ��+���ҏ����� ��,�P�b�t������� 9�Ο�����(��� L�^�p�������5��� ܯ� ��$�6�ůZ� l�~�������C�ؿ� ��� �2��_�_h�o ���o����������� 	��-ߛ�9�c�u߈� �߽߫����ߣ�*� <�N�`�r��Ͽ��� ���������&�8�J� \�n������������ ������4FXj |������ �0BTfx� �+����// �>/P/b/t/�/�/G� Y��/}��/Y���?'? 9?K?]?p?�?�??�? �?�?�? OO#O5OGO 	�~O�O�O�O�O�O�O 5/_ _2_D_V_h_�O �_�_�_�_�_�_u_
o o.o@oRodovoo�o �o�o�o�o�o�o* <N`r��� �����&�8�J� \�n��������ȏڏ ����/�/4��/X��? ]O{�������ß՟� ��g��/�A�S�e�x� ������oO����� ,�>���P�t������� ��ο]����(�:� L�ۿpςϔϦϸ��� Y��� ��$�6�H�Z� ��~ߐߢߴ�����g� ��� �2�D�V���h� ����������u�
���.�@�R�d�� ��*default�q�B�*level8˯%�ï������� tpst[�1]��#y(t?pio[23*� u(������	�menu7.gi5f�
�13�	��5�
��
�4	u6�
گOas�� ������//'/ �K/]/o/�/�/�/�/~F"prim=��page,74,1�/�/??)?;?F"��&class,13@?v?�?�?�?�?M?_25�?�?OO0OBOE#T<�?|O�O�O0�O�O�/�"18�/_@_%_7_I_TO^26P_��_�_�_�_�_��$�UI_USERV?IEW 1"�"��R 
���_N�oo�m8oaoso�o�o�oLo �o�o�o�o9K ]o�,o���$ ���#�5��Y�k� }�������V�׏��� ���,�>�P��� ������ӟv���	�� -�?��c�u������� V�`�ʯܯN� �)�;� M�_�q��������˿ ݿ����%�7�I��� V�h�z�쿵������� �Ϡ�!�3�E�W�i�{� ߟ߱������ߒ��� ���S�e�w��� >�����������+� =�O�a�s��(����� �����'9�� ]o���H�� ����0B� }����h�� //1/C/�g/y/�/ �/�/Z�/�/�/R/? -???Q?c??�?�?�? �?�?r?�?OO)O;O �/�?ZOlO�?�O�O�O �O�O_�O%_7_I_[_ m__�_�_�_�_�_|X