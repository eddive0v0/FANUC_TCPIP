��  �A��*SYST�EM*��V8.3�0340 11�/9/2020 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  �  �ALRM_�RECOV� � � ALM"EN5B��&ON&! �MDG/ 0 �$DEBUG1PAI"dR$3AO� �TYPE �9!_�IF� ` �$ENABL@�$L� P d�#Uژ%Kx!MA�$iLI"�
� OG��f �%CAUSOd�!PPINFOE�Q/ �L A� �!�%/ H� �'�)EQU�IP 20N�AMr �72_O�VR�$VER�SI3 ��!COU�PLED� $�!PP_� CES)0s!o81s!Z3> ��! � $�SOFT�T_I�D{2TOTAL_�EQs $�0�0N�O�2U SPI_I�NDE]�5X{2S�CREEN_84no2SIGU0o?|�;�0PK_FI� �	$THKY�-GPANE�4 ~� DUMMY1d�TDd!_E4\A!R��!R�	 � �$TIT�!$I��N �Dd�Dd �DTs@�D5�F6�F7�F8�F9�G0�G�GZA��E�GrA�E�G1�G1
�G1�G1�G �@!�SBN_CF>"
� 8F CNV_J� ; �"�!_CMN�T�$FLAGyS]�CHEC��8 � ELLSET�UP � $�HOC0IO@� }%�SMACRO�ROREPR�X� D+`�0��R{�UHM�P�MN�B�! UT�OBACKU��0 �)DE7VIC�CTI:0�A� �0�#�/`B�S�$INTERVA�LO#ISP_UN9I�o`_DO^f7��iFR_F�0AI�NA���1+c�C�_WA�d'a�jOF�F__0N�DEL��hL� _aAqQbc?Yap.C?�Y`�A-E��#%sATB��d��AW{pT $DB� g"� =S�$MO�0B x!kq� \� ;VE~a$FN!�p�d�_�t�rdTM�P1_F�u2�w1�_~c�r~b���MO<� �cE D [�mp�a���REV��BIL0�!XI�� �R  �� OD�PT�$NOnPM��I�b�/"_�� m�蘁H��0DpS �p E RD_E�L�cq$FSSB�n&$CHKBD_YS�r�aAG G�"$SLOT_�H�2��� Vt�%��x�3 +a_EDIm   � �"���PS�`84%$�EP�1�1$OP��0�2qc�_OK8ʂ� e0P_C� c��+dR�U �PLACI4!�Q���( �a�p9M� <0$D������0pB�UOgB,�IG�ALLOW� �(K�"82�0VAaR��@�2�sBL�0;OU7� ,yq�`�7��PS�`�0M_Ox]d���CF��7 X0GR`0�z�M]qNFLI�<���0UIRE��$ށwITCH�sAX�_N�PSs"CF_�LIM�t=�SPEED�!���P��p�PJdV���u�u�3z`�P6��ELBOF� �W��W�pH� ���3P�� FB ���1��r1���G� �� WARNM�`d܁�P����NST� CORz-PbFLTR۵/TRAT�PT `� $ACCQa�N �r�pI�o"���RT�P_S�r C�HG@I�Z�T(���1�IE�T�Y1�݀�� x pi#�Qʂ�HDRBQJ; #C��2��3��U4��5��6��7��U8��9s!�k�M$��	3 @F TR�Q��$�V����C�FN�_U�pY�k�OpT <F �������#�I2q�LLEC7�>"MULTI�b�"��A!cj DET_��R  4F S�TY�"b�=*�)�2��o���pT �|� �&$L�>�+�0�P��u�!TO���E`�EXT�יၑ8B���"2����
�t k0F�RLƯ�r�q���� !D" �M��Qm� �蠋ck�����"��G�1�ց�qM���P��! �����# L0	����P �pA��$JO�B,�ǰR�0�TRIG��$ d��������� �K� l��弧�o�_M�0b% t2��F� CNG0A�qBA� ��x��
�!�v��� ��z�0�P�{`�R·&ΰ@f�Pt�a�!��"J!�S_R��rCJ$�T(J)�D�%CH ӽ��z@h�P�Z�@ '.�RO`�&��סIT�c�NOM	_�`���S ��pT(�@�݉��P�ǭ��RA�0�2x&"�>�
$TFV .w�MD3�T���`QUC1[�g�'�Hgb
�s1q*E���\Ѕs��qŦgAŦsA�YN�T�q�P|pDEF2�!)��G�PU8/@0�����AX��Ģ��eTAI~cBUF�ņ�|psQ* � ��'�PI�)*�P\7M[8Mh9� �k6F\7SIMQS�)@KEE�3PATѠ"�%"�"$#�"��L64FIXsQ+3 ԭ�AdC_v���1�23�CCIh��5�PCH�P�2ADD �6,AE,AG,A!H�_�0�0_,@�foA )�ԀzFK� '�=$#�"t��4E��, l����7zpF�CE�C!F +HS�EDIS�G�3��-�P��MARG8���r%�FAC
��rSLEW<���xX;�M��MCY.����pJB����
aC��Wv��U�W/ ��?�CHNS_E;MP��$GE gB݀_} ����pP�|!TC9f��y#a��� NdW#%I��r<��<��JR�И�SEGF�RoPIOj�ST�`�LIN׃�cPV����!�$0�����b�'��b�B��1` +`��	��a	` k�a�Pܠ��At��Py�QSIZ���ltKv�TVsE pz�y�aRS %Ѽ�uc@Q{k�|�`�x�Z`�`Ld�| `�vCRCɥ��!����t�`�%�9a˭9blMIN@Q�9a7��q�D�YCk�Cz��le��50��p ��EV���F*ˁ_leF��N���P�Q۶�X%+4,���#0|!VSCA$�} AY��c1G"�2 �>�
/Ψ`_rU @�+�w][��i %�7���R��3� ��ߒ߱���5ġRޟHANC��$L�G���*1$�0NYD�סAR�0NK`�a�q��acm�ME�10��n�A0h�RA��m�CAZ����X%O`�FCT���7`�v�S�P
ADI�O ���u��pWP ���������Gv�B�MP�d�p�D&ah�AcESf@̓�W_P��BASk�s��4 � �I�T�C�SX@�w�5��	-$�1�T��?s�Cb�Ny`lBP_H�EIGH71��WI�D�0lVT�AC��u�!AQP0� �\��EXP+�L�@��C}U�0MMENU���6��TIT�1�	�%��aǱA1ERsRL���7 \��̉q��OR�D��_I�DG��QUN_O|d�L $SYS����4�ő�Iϡ	�E�VG#�a��BPXW�O����8��$S�K�*2���T(�T�RL��9 �� AqC`�u䈠IND� �DJ�4 _Z�*1XK�*�W�PL�A�R#WA.�tТSD�A���!�r@Y�UMM3Y9�ª�10����d���:	�A1PR�qw 
��POSr���; ��[$�$�q�PL��<��ߪS@��=�'�Cr�>4�'�ENE�@�T{�?S�S��R�ECOR.�@H� �O�@;$L��<$��62����0�`_q���_D9�W0ROx@�T[���.�F��������P�Ac���bETURYN�V�MR��U� v��CR��EWM�b�mAGNAL� 72$�LA�e��=$=P�>$P٠= #?y�A<�C���@�DO�`����:�>��GO_AW ��MO�a)�o���C�SS_CNSTCY�@A L� ^�C`L' ID[^�2
2N��O����ـI�� B P�NPRB^rzCPI�POvI_BYȀR}�T�r��HN{DG.�C H��DQkSP�s*�SBLIO�F��0��LS�D��0N0�	3FB��FE���C��жE�DO&a-sO�MC`{P�4�C�rH��WFP8B���SLA�P�F�bIN� �N3����G� $$���P]��v��v�ޕ���!o�"��#CID�&L�&W�"�;$NTV*3"VE 4��SKI��as$�3�'2�&aJ�&a<M�mdSAFE,d�'�_SV��EXCL�U7ѻ���ONL`�#YcL���4���I_V8���PPLYy�R��H[0'3�_M@�NPVRF�Y_S�2MS�O@��k6�1�~3�#�Ot !5LS�E��3�5�£1�`%�P���$��t5�%� 3Hy��TA2�DPι� �Q�SG�� I � 
$CURB�_�
�B �������#H��3F��UNM��DZD@���l�{IxA��J��F	BEF��IM�J� @F]Bk��pOTb�k�ԋѭ5�׿P��и@M� NI��K���
RwPA!(TD{AY��LOADj��R�ӵ2 �EFV/�XILy��q�}�OhPe�D�_RT;RQ�QM DF�����P�r�S`�ThU 2L�`���Qk�P8���Q�QN 0�A�QaA�t�R���DUb���"�CAB�aO��B�NS�QW`ID��`PW���U/q� V�jV_�P�P���D�IAG�1�aP�O 1$Vb�HuTl�@�u�t� �j���rRp�lDQ�tVE��Y@SW�ad�p7`U2�PM�p�QOH�U�Q3PP�`�sIR���rB��Fb�S��q��q�@ 3r��-x ��-uj#e��PO��P���uRQ�DWuMS���uA��u�b�tLIFE Z��C�p���rN�q�r��uxA�s�rI�xBCVp���NC�Y����FLAW�y@OV����vHE'ArSU'PPO2���rS�1_E�)E�_Xf�h���s�Zp�Wp�p�s�0��xA���XZ����V�qY2ˈC
�T��D���eN됕exAJ� v_��q�/����Q `[ CACH9E��3�SIZ�v*���"j�N� UFFIo� �p���Ե3���6��dat�D�M����R 8�@K�EYIMAG*�TM�ᄣ��D����>��OCVIE�`�'S ���Ll$@)#?� 	��%����T�P�ST� !��`!��@!�VP!�|�0!�EMAILy��1Q��� _FAU�L��U� �9��C�OUz ��T��|aV�< $��zS��PC`IT�#BUF@F�)!F�Oy�o�D�	B��nC($�������SAV�Ţ�`� ��`���|FP
�z���d� _���"P_�#OT�����P[0���� B��AX��-�I����Wc7�_G�s��YSN_$q'�W�RDuTY��#rMb�T��F�fP^@D�&�X������g�C_��&�K��8�4B�3��R��2�q��D�SP���PCy�I�M�pÖ��#�Æ`U`M�:���K0d�IPm#0�q	�o�TH��=�c�mPT��p�HSD=Im�ABSCz$��o�V� �Я�&�`��QNV�!GO�&ԑ�$mƸ�F�aаdR������SCxbk(�M�ER4�FBCM�P3�ET�1�Y6��FUX�DU���\���%2CDf���z��u��R_NOAU]T�  Z�P4 ��"U�IUPS�C�א�C�1ϱc�㍰��[H *�L t�3���� �@�0�#�����A��@VQ��1�扑��7��8��9���p���1���1��1��1��1���1��1��1 �2R�2���2��2��U2��2��2��2��U2 �3�3��3��B��3��2����3��U3��3 �4�_�sXT�aQ\ < ���I簉���3�FDRxd]T��V�0���r�.�rREM�`F��r�OVMI�>AGT7ROVGDT�gMXvING�fNuaIND��r
�<�а$DG��:s�p��u�aD�VpR�IV���rGEA-RI�IO�eK7�tN�%(hQ�x0h `�>�sZ_MCMÀ�q�;�UR��^ ,<�1? �� s?� �a?�!�E�0�!	A����_�dP}pP���`RI��դ$�aUP2_ g` VPģTD��@�3�#?@�!�'�%�%wBACܲa T�hŢڠ�A);@OG.5�%�CT����IFI�q���x�:pC5PT�V��FMR2
bO �3LI��3#/5/G/P^|��u7_��"�R_�A�԰`M�/�-DGCLFuD7GDY_HLD�!�A5�v��tz3�c�P��9 T�FS]��d P� �B�0|��а$EX_�A��H�A1kPl���@3�[5V�G:�
e� ����SW�O>�vDEBUG4WR��eGR� �U��B�KU��O1a� pPO�P�YoP��lBUoPMS�0OO���QSM�0E��!��� _E f �Ő �TER�M�Ug�U���OR�Ie0�Qh�W �S�M_80Ţ�Pi�UV_F �TAiji�UP�k� -���f$�Ua`g�$SEGfjx@EL�TOV�$USE.��NFI"��bn ��q+�d]dh$UFR02���a���	@3OT�gU�TA ���cNST`PATx��?��bPTHJ ����E�:��АbAR�T+��e|�+�V��aR�EL<z9�SHFTp�a q.x_SHI�M^���f $`�x9j)A�0OVR��ǲ�SHI_p&DU4� %�AYLO��Aֱ�I�ѻ# qk�%�k�ERV���q�yz��g�`<r4_0&���_0RyC�!9�ASYM	��9��aWJ�g��E �#*qV���aUz�` ֱ.u|���DuP���p,YѪvOR`M�3Z�GR�Q1Tl�oR�V��`�`AؐB��m ��>�b671TOCb�a�QT!k�OPZ2����}���303O,YߠREM�Rm�9��Oѐ$�reT�R��e��h�Fq/4e$P�WR�IM���rR9_C�#tVIS`sfb�UD�#fsSVW��B��b n� $�H.56�_ADDR
�H�QGr2�'� ��t�R��~�o H� S��Q�4_���0_���_���SE�A¿��HS��M�N�Ap `T���_����OL����v���ּPACR�O���aS�ND_C�����qٔZ�ROUIP���_X���@��1��25���?�4  ?�<@���?���?���6�2AC�IO��W��D:���J����1Sgq $� ;�_D� x�PM���PRM_.��H��HTTP_��HQar (�O�BJE��"�/4$��LE�c��s� � ���AB%_�T�SS�S� ��DBGLV��KR�LÙHITCOU��BG��LOF�R�TEM�ī�xe��a7f�SSQ ��JQ�UERY_FLA����HW��aQat2Z���F�PU���IO�h����u�����ѿ� �IOLUN2u��
@C���$SL�2$I�NPUT_�1$ă�i�P m�D�SL��Qav��gߢԝ�=��s�=��IO�F_�AS�Bw%0$L :0'�:1�q��U`|p§aTժ�_��pHY�� �������UOP�Ex `��>��� ��hᣐP�Ã��^����x�.� U}J	y � � ;NE�wJOG�g��7DIS�3J7���+J8��7!PI�a��>�7_LAB�a3�x�����APHI� �Q��9�D�@J7�J�� �@_KEY�� �K�L�MONQaz� $�XR����WAT�CH_� �s98��E�LD.5y� n�E{� ��aV�(���C�TR@s����%R� LG�|���~DSLG_SIZM��� &�@%��%FD0I$;�Q2#�P =/" _�+��@���ЩR ��P��S���� �ťV" ZIP�DU�r��N��3R}J���@P�A��]�"d0U�-�L6,7DAUREA��/�h^GH0��!���BOO2~� C��ӐIT�Ü>@���REC�SCR�N����D����'�MARG�2Ҡ����ӐN�"����S3���Wp���A��JGMG'�MNCH����FNtd�J&Kp'PRGn)�UF|(�p|(FWDv|(HL�)STP|*�V|(e0|(�|(RS"�)H�+��C�t�# y���1P#'G9U籐$@"'�r0&���"G`)�WpPO�7�*��#M�07FOCwP(EX.��TUIn%I�  #�2,#C8#Cl p!��p��v3@���p�N�sANA�҉b�p�VAI��CLE�AR�vDCS_H�I\T�Bu��BO�HO&�GSI�G�HS�H(IGN; ��Mm!���T٤�@DE�(4L1L\�C���BU�PR`����pT4B$F1EM������rRQa����pW��\Ρ4�OS1zU2zU�3zQ�_�AR`� ����΁�esԲsԗIDX�P�r��O��P��a�VST?�R�iY��a �$EfCkW��&fp9f�V��V�� L�� �_�#�|p��U���ו�E��֕YU�_ � �� .������c �MC �{ ���CLDP?�>J�TRQLI�[�8���i�dFLG���`���srAD��w��LqDutuORG�� !21r��vyxu��t���dд� ���t"5�du� PT�`��bp��t�vRCLMC��t}��y����MI������ d)�QR�Q����DSTB�P��P [��h�A�X�bi�k���EXC+ESy�;�M��U��O��ddat�=��V��Z�]�_�AW�\��������`K�B� \�����$�MB��LI�I�R�EQUIRE�cM�ON�
�a�DEBU���EN�ML�`MA� ڰ ᛐ�����q;�ND>S���'��ړDC��2:IN�7RSM�����@N���F3���ҁȑPST� �� 4}�LOCf�VRI���UEX\��ANG�RY�;�ODkAQA�K�$t�1RBMF��]���Y��b0�eǥC�SU�P�eJ��FXS�I�GG� � � ���b�wÓc:6�d���%c�?��?�.�<��DATACWk�EE��E�����N"R�� t��MD��I��)���@��-���H�p��ᥴX�!�AN�SW!��`Q�1��D���)|��� ��� -ÀCU; V� pLx���LOj�����$5�W�3�E���UƼMê�MRR2B��O� (E�NA�q� d$CALI�a��GvA��29�RsIN� ��<$R���SW0���)�AB�C��D_J2SE�u�Y���_J3��
���1SP���Y�P����3�"��Y�BJ�J�CZ՞r�O!Q�IM��(�CSKP z��1oC��Jq(��Q�ܺՠպհ�e�_cAZ�rV���ELQ<U��OCMPs�)�����RT��G�11���5��P1�9�f�:G�ZE�SMG0}�L�Օ`ER�����PaA �S(���DI�v)�JG�`SCL��n��VEL�aIN�b@��_BL�@Y��䄀�Z�J��������p�x�IN�ACcR�@��	"x��f`_u�!�<���<�܂�F���x�DH��;����iP$V����'A$d�b��P`���qy�B��H �$BEL��|��_ACCE�� x�����IRC_�����ppNT�Q�S�$PS���bL   ��&s�	1w@
PATH��_��_3..���_wQ�� Ȗ�rb�CC ��_M=G !$DD���`�FWE�~����������DE�PPA�BN6ROTSPEE�{Q�`��{Q�DEFb���. $OUSE_��BCP���C�0BCY���q s�YNA�A�}y�ܼ�}MOU�NG�RR� O��Q�INC�m���h����i�ENCS��d�Y��&��f�# IN�RI0.%���NT����?NT23_U��`�^A#LOWL�A~0��`�a&Da0Y�C����`���C,�(&M3OS�@�MO�ǀ��wPERCH  ~#OV�� �'�Q�# F�d"&�F��
�gm $�@w�A. 5LADwӀ�v�)%�d*_6z&T3RK���QAYI�3 쁏1.�5�3n������PMOM Bh�� sp"�W�����3a�zR��DUЋS_�BCKLSH_C .!E��&� �-�?D��JJ���CLAL�BP'"�q�0܀|ECH�K�`�US�RTY�J�N����T:Seq}�_�c�$_UM���IC��C����C(LMT�_Lwp� ṮWE]&P[P!U�,�5A�+0gT8PC��!8H�`|���EC��p�bXT���CN�_��N���V�SF���)Vg�a	'|�Q�.
e�XCAT�NSH������eq
A
&`F�/F�Z� PA�D&�_P�E�3_�`����6� �a�3�d�EJG0�p���cO OG�W��TORQUY/Ւ#��9� ?��"��� r_W�5�4C��<t��;uT��;uIC{IQ{I��F��.qaҐxpѽ VEC��0b�Z��r1�~p���s��uJRK�|X�r�v�DB��M��:�M�_DL��:2GRVBt;���;����H_L��b i�CcOSv��v�LN�p �������d���mq׊Ō�q�Z���&�cMY�����TH���6�THET0j%N�K23��`��㣀C�Be�CB��C��AS���mt����e��SB��p�GTS��(C�m�=�cM�<�ԃ$DU�@C7 ����� ���QF�s�'$NE��ؠI���C)���T�AX�����8h�s�s�LPHv�_�9%_�S�ңŅңԅ@_��������V��QV����VʪV׫UV�V�V�V�V�H��E�²��?aTٸ׫H�H�H�UH�H�O��O���ONɹ�OʪO׫O��O�O�O�O�F_�����Ņ�Ė��SPBALANC�EQԃQLE͐H_X�SP�9�ņ9�>ԆPFULC=�dҰL�d�ԅ&�1��U�TO_�@�eT1T2����2N�A��? �Ԗ��1f�D�5���1�TP0O����,pIN�SEG��!REV8�փ "!DIFy5K��1�0��1� O!B&�lAE��72p?��A$�LCHWAR���AB�a�5$MECH��%�����FAX�1PJT��z���З 
��q�n%ROB� CR.���R[�MSK_|���� P ��_WR��r0�?{41	b4 20�1#JD0����IN��MT�COM_C�p��  � 8��$NORE$#����t���� 4�0G�Rr��FLA�$XYZ_DA���nC DEBU�� X��t�� 0�$uwCOD[A ����2���0$BU_FINDX2��C MOR#�� H-��0���FB �0�8JD$����QV6PTAAp+�2�G6� � $SIMUL�` 1x3�3OBJE;�>�ADJUS�� OAY_I�A	8D��OUT�`���0�_[FI�=@T+p 4 ��X�3p�3�A�5DrFRI4(CXT8ERO�` �E3q[0�OPWO��p'�, SY�SBUq�( $SO!P��A�U�3��PRUNv��PABC�D���0_� NR�X�AB��PP� /IMAG[A-�G��P�IMY"$IN�,��!#RGOVR!DM�� �P   #`W�L_��an%�B��PRB5PX�`QMOC_ED/ �� PP�Nq�M�"OQ@MYc19NQ�M!SL;��'� x $OwVSL��SDI{DEX�S�&�SP1�"	V3p�%N1q�0�378�"A�$_�SETp'� @0�0K2��AARI�� �
^6_��j7�1v1p�5� �P �<yT���`ATUS@$TRCI�H%N�3BTM�7�1I�²$4NQ�3� '� �D-�E��"�2z�E�v��1!0l@�1EXE�0�A�!B*B�4S31�Z0.��0UP��9As$Y�' XNN�7�q�$�q�9 �PG���� $S�UB�1��1�1�3J_MPWAI,`P	3��ELOP����$RCVFAIL#_CH��AR-�����Q�P�T�U�R�_PL�3DBTB8�a�R�BWDV��3UM�`TIG�( ��4`TNL(`TjRARm���`
p	1XQ¬ E�S�T�R�ADE�FSP�� � L-���P_�P��S�UNI#�7�PmARX1@��3�_L�P�1F2Pw�&����`�� "<0��)ОNU�K�ETb(p��`P�^R&� h� ARSIZE� ��1���naS� OR�3FO�RMAT��TTCOX� ja�EM���d��SUX�2bLI�OR&�  $>��P_SWIu�����fLLB&��� $BA�`1�ON9AKPAM�0=y��BAJ5���2r�68v��_KNOWH8cNrA�U9AߐDx�� �PDC�ryPAY��[�t���y��wZ�sL�1���PLC�L_$� ! A�s,qv�tb"�v=F�yCRPO�z�2&�tES���wR4��w��tBASE$�JL��W�_J�qK�mA��fBu��r�qG1�MAX4P�`AL_ � $�Qh 1qT�!��C[�D�sEfr��J3����� T� PDCK� ��CO_J3�������
�hr���� ���C�_YQ�  � �\� �D_1�z2�tD���n�^���m�|�TIA4��5��6[�MOMS ��ȓ��hȓ��B�@AD��p억��PUB{AR͔����;�e�#��` I$PI�$�QM�=q�wk�B1��yk���������iqR�M�q�!Ħ~AĦ�A�
��9d5SPEED�G�b��E�T� �T�EP-�C��Q8+�Q�ESAM(�E������Ep{� m�$�� k�~@ Ƕ�P_�ֹm�k�v{���ŵ��,H��ǳIN̚�c��1���B��W�.�W�w�GAM�M��1��$GE�T9" �D;�u
���LIBRcA�RI.��$HIb@_=!�0$k���Eh ��A����LW��4�+��X� �7���wP��CEUv�[ �0 �I_b�xu��L��������ȓu��ٞ� ��$Ј 1�*��I�0R��D\��kAT��LEf�=q�1�M�7�ୄPMSW�FLTM��SCRsH7�����!��~B�d;SV&�P� A ������#S_SA�qs$��eCNO;�C �1fB<�����K��� ��S�C���hrǥ��m�D� a���� ���в �����C�����L���s ��`MJ�߰ � ��YL(i�K���^SJ�| v!6O�K���BK��- ��OW�� �9���M$P���p����Dc�"��1�~B�`M��T2� �� $-�$$W� �%ANG"�q�  ����!��5P�&��o����c�#��X`O"���Zz�`�@n� �y�OM��+�(�:�L�^�p����CON@�eL;�_�B� |ၰ��ș @&��@&�࡚m'X&8��.��� '�⥴�`X$$Pma��PM0QU�� �� 8#`QCOU����QTHYPHO�/� HYS�`ES�-r� UE� ��S`O��d�   $P��@�Ŋ2UN�0br�@O��  � P�p�45�E��C�RROGSRA�1A2DO4�45IT�Ё1F0IN;FO�� %0g;��1AȬ!OI�2�{ (�SLEQ�� �1��0k6E1S�НD�� 4#`ENA�B"20PTION��C�T̢/G�TCGC]FA� @#`J$P���<2���RdH00OBGb\�ED�@  '� �{K�q�35��E)�NU�G�H�AUT�ECOPAY�qI0�L���M���N�@�K��PRUTj �BNV@OU�b�$G92DTH�!R�GADJ��bbX_ �R$`pV�
pVWnXPnX[�pV��`Pz�N��_CYCZ"ZSNSE�$ ΂�LGO���NY�Q_FREQ0�W b��a�d23L�p�b��PnQÓb��5CRE����#��IF��s3NmA��%?d_G��STATU' ��*7OMAIL��YsIN��$LAST�a���T�ELEMA� �|��GFEASIA ����H �b�1���f;B����I�0���R=q0�!� R�rAB+A��	Ex0�V�a7vW�Cy���1�U8�I0�p�d�lvRMS_TR s��@��sr7�z��a�ktB�R�/ 	~�b 2� =� _+��ve��w�r� ��fe��c�G�DOUda3;�NHC�RPR	 z@��2GRID�1�+CBARS��TY�C�ROTO㐾����&0_[d!�P��B��OxD� � �0�PORa3��[�.��SRV_`)˄ÆDI�T^���������4��5��6J��7��8ぬ!F���A�#0$VAL�URs���d�q_�D�� E��u1��1aa��=@AN�㉒�qaR�@a��TOTcAL��1��PW�S�IJ���REGEN����#XxxI3e%!���� TR^s0���_!S��^���CVnQ�D��B8rE�cN��!��42�@ÓV_Hk�DqA�~���S_Y
�rfS��AR�2�� <RIG_S!E�ch�Â�e_80���C_v�`�ENHA{NC�!� p�q�Eqb�ý�INT���� F.3MAsSK��ipOVR�#P� N��`a
�_�*6^�M��B[��f8���SLG����� \ ��eH ���YSq�dDE�U�� *7Ő�%��U�!��TEj  � (7��҆�J϶�"cIL_M!d��P㈠�TQ� �Ë1rpj�jeV��C��P_���op��M��V1��VU1��2�2��3�3��4�4���ᄠ��������s��IN��VIB� �İ����2��2��3��3
��4��4�ؾ���#" �������%��׌ՠ�v��PLv`TOR� ��INb�����  ��p��MC_F,� 	���L����B�ڐM�IB���#�� 1 �)���K�EEP_HNADED��!��<p��C��_`�䂁��H ��O �!��P������G���REM���쑥��;�R�W�U[de��HPWD  ��SBMo���G�1��2�� H COLLABu��a�����h�ؑEb�0IT��p��0��� ,� �FLbq$SY�N��M�C��~d�UP_DLY�=�#2DELAJ ��nbY� AD�;�� QSKIP�� Ļ�60ODD���t P_60_2�g0^  ����		Q�	��	 %��
2��
?��
L��
�Y��
9�Q�J2RT�P��CX]pT�SY��X]P��Y�1��� RDC��b��K ��@ReCg�R4ape��"d��RGEr@8sl�:�FLG�!P�a�SW�I��SPC��3�QUM_Yt�2/TH2N&�# L� 1� �E�F�@11�!� l������C��AT 4�ET1��7s"k0o4j!�@Y�j!<3\�HOMQE�"�P<$2D"�J/@\/n/�/�/�/�'3D"��/�/�/�/?!?�'4D"�D?V?h?z?�?�?�'5D"��?�?�?P�?	OO�'6D"�>O@PObOtO�O�O�'7D"ֻO�O�O�O__�'8D"�8_J_\_n_�_��_�%S��1�9 ��q=#$���S�E��ٷ��Lbݖ&JcIOq�jiI�P���GbPOWE��G� 4` wGb�ה ��b$D;SB�GNABqՔ�E C) ����S2;32Pe� ���Uy�P�ICEUQr�t�E3 ��PARI9TáՑOPB��oFLOW�TR`��c�3���CU+pM���UXTn���U�EORFACtC�Uѐ{pRSCH�q'� t����_p�f�$����OM۠�9�A�T>���UP%D�A#�`T+`҃�*�� �x�s!��FqA������RSPqp�Q��� !�X$USA ���Y�EXmpIO6��pU�	YE��b_�ª�B�#qF`�WRp��_�YD������VFRIEN�D���UFRAM�δ��TOOLȆM�YH����LENG�TH_VTE��Ix���[�$SE�`~��UFINV_�@��5aRGI��N�ITI���XX�l	�J�G2J�G1T� U�D�d�u���_Â#O_p�py�ၻ��"n�C	�zŔ�C ���ʖ �G��zr2�� @ 9�qC����d�wu��ysF� ����p��X n#�E_M�pCT^��H��f��<u6�	�G�#WV�z�G���Dh LOCK~�U� �������$� �2���~�D ��1T���2��2�3��3���:����V��VP=�"�=�F�V��!Р��/������p� xṿ����Prƻ���������E����؅�!��AC�PRs�!�}�S���`��K�r
��a� 0 5�ؠ�V��ؠA���	������
MŽS��� ح�R��qda��$RUNMN�`AX2q��A���L�+"��THIC�x� w �u��FEgRENg���IF���x���I����V��G�1&�*Ԅ�1ٲ[�nI�_JFR�PR���
��RV_DATA�q� RD�[- 
�AL� �x�Α �b{�  ?2� �S��`?�	� �$ Z="GROU��!�TOT����DSP>��JOGLIYs�'E_P�PrO��\�7`��bvK�p_MI�R�.䎐MQ�O�A	Pp��E<�o��t���SYSE�ib��PG���BRK���v$ A;XIa  �⃃����Ҽ�A����H�B'SOC��T�N���{16�$SV1��DE_OPNsSFSPD_OVR4 ʓ���D� �OR$+��PN�P,�F��,�6�OV�SFa���d�$�F}�ja2㒓���ҁibLCHH\R�ECOV�n��WbE�M����RONs����_���� @��9�VER��n�O�FS9�C�Я�WD�E���A����Rh��T�RBq6aY�E_F�DOh�MB_CM4kS B��BL��.�u��8�V摁��p�d��]�Gv��AM��`i ������_M� �[r�ec T$CA���D��HB�K�q�vIO��8,�a��PPA L�1\D��bDVC_DB<���q�b���ja�1���y3���ATIOi`jqcp�U�� �efCAB�����J��������__p�vS�UBCPUP�S v��`_��p"�`'}����b"�$HW_AC� Ip���'ɣAx�~���$UNIT���� � ATTRIx���"�CYCL���NECA�Y�FLTR_2_FI#�0�h��f��LP$����_SCT��F_Ʋ'F_�,E2�*FS8�a��"CHA��-7p�1�Pr�2RSD  `�b����Q�`_T��PRO�MFpEM�	`_���Ts2��c s2���5DI&�~�tRAILAC���M��LO�����5��������P�R�S̑{�dAC�p	��FUNC!��RIN됫�|��@�DEqRA�@�� ��C7`�CWARB�	BLƑ�G�DaA�K�!�H�HDA��0�AX�C�ELD�p𐒡@S���A�@STaI��`U�ѓ�$<�gRIA�q�bAFQ P�a�S��U �����3MOI� PD�F_ꀔ��qHpLM��FAE�HRDY.]�ORGEPH�0���|� P�UMULSEP���`'���0J(��JC�X�S�FAN_�ALMLVBs_aW{RNfeHARD����v�䐟p�@2$SHADOW��0��a@�b��_`+q�ї�_���vAU�Rx4\rTO_SBR��e����j� ��A	sMPINF���!t6Q'sgREG���aDGBPb��V�p.�l�FL�%!���DAՀ_��P�CM��N�YƧB �V  ��� �]���$N�$�Z�� �Ҭ����7� �|�EG���ӌ��qAR��#��2p?��wP��AXE��wROB��RED���WD���_F���SYм�!���h�Sr�WRqIE��v� STR��(�`��7�E�!�����a��B����@C]D� OTO7q����ARY����.A�̟�#�FI��9�$�LINK�Q���Ry�_���6��N8�XYZ�bB�7P�'OFF
 �7�+�%�B��yB�����0}@��FI� ����h��yB
�_Jဓ�5�����`Ȅҋ8���H�TB�b�CL0x�DU �9AETURa`XgSW���brX���FLz�@��#�pu�Y���3\���� 1��K�M����31�DB`%8��`'2ORQ�6�� �C��}�DB��>��P���%�����\q:�OVEA���M90=ѻs[��s [��rZ��`X��aY��  X�O�~@91�P��B�F� ���=�S�B�_���s�����ER�A	BEBE��� QC"�Aб�����E�2��Q&QAX���Q� �! �|�A��+a����� @@��O���n������N���1����`��` ��`��`��`��` ��`��`��`�!���� �Rg�DEBU�#$�A�c�2���3�ABGE�;�V�" 
�Ҷ�� �z!$�
�$��$�@A $�O�$�n�$��$�N���T#��R����LAB⬒�� �GROh0��l� B_�1 	ƞ�>��`����8���a	�ANDàE @��<���aF� ���q��Z�Qi�� ;�NTq`�cR�C�1=���
�� �pERsVE���p� $q�ڱ@A�a!��PO �`X �����Q�p��p$��TREQm�
��Q����ƑR2�oP@_ �� l=���fESRRҒ�IV�����gTOQ����L�%��Ď�z�0G��%�%�"��?�!P � ,��2 뺱R�A� 2� d��D�p�  ��p$O��2�Pvµ�OCQ� �  }YCOUNT����FZN_CFG���� 4� ^v2T��d�"���m W k!�E�s� ��M �08b�����X��0�CFA~P���V�XA�@�����0���O rA�P�b�pHELkp~N� 5ސ�B_BAS�#RS)R]vm@;�S�!YQRB 1�B 2e*3e*U4e*5e*6e*7e*98�5!ROOGP� ��:�NL�q)�AB���@C ACK�I%NT80�sU�``x1�)_PUA��b�2OU��P�@^x"#��y0��b�TPFWD�_KARlfpZR�E���PP�&Q�@QUE]zROB�2����`�aIb`�"#8�$C80Bv8�SEMա�6t�`A�STY43SO�0�dDI1�@pr�1aǿQ_TM�s�MANRQAF8�E�ND�d$KEY?SWITCHS3h1�#A�4HE2�BEA�TM�cPE�pLEPks1���HUg3F�4�h2S(DDO_HOeM�PO�a� EF"�PR���rS����v�@�OaX �OV_Mx���`pPIOCM$���7���!%HK�q� D5�_w�	U�b�2M�p�44�%��FORCcsWAR��R9�##OM�p �� @��˓�`U���P�1�V2�V3J�V4��Ox0�L�R��^xUNLiO.0�ddED�a�  �$$CL�ASS `���4.a-�-� #`�S�0+h9`;��?aIRT?�,o�>`AAVM��K �2 je� 0  �5�5a�o�h�o�m �l	�m-�Bk`��o2v7u�l V}b�ah���t{`sBS4�� 1Li� <� �� �2�D�V�h�z� ������ԏ���
� �.�@�R�d�v����� ����П�����*� <�N�`�r��������� ̯ޯ���&�8�J� \�n���������ȿڿ������rC`�AXؙ� `���s  ��%�IN.�@�$�P-R�0XEQ�}�`�'_UPMIl�ja{`9L�PR ji`���tLMDG �g�`��PIF �k`d��0� B�T�b�߅ߗߩ߻���, 
���n� �o�0�B�T�g�x��������yNGTO�L  �{�pA �  ��
�{`Pd�O7 �� ��=�O�a�s�6b� ��u� ��2b�������������&J4Z���� �������*<N`r��zP�PLICA�1 ?�je}�����Handlin�gTool � �
V8.30P�/58��
8�8340��F0!�755���>�7DC3������ޝ��FRA� 6�*-  !�� TIQVqŵ>��#UP�n1 ��\�PAPGAPONf`�.za� �OUPLED 1�i� /03?E?�W?�_CUREQ7 1�k  P�a7a<�n�?�d}��3�3b9b ���4H�522�:HTTHKY�? Kx�?�?ZO�?6OHOfO lO~O�O�O�O�O�O�O �OV_ _2_D_b_h_z_ �_�_�_�_�_�_�_Ro o.o@o^odovo�o�o �o�o�o�o�oN* <Z`r���� ���J��&�8�V� \�n���������ȏڏ �F��"�4�R�X�j� |�������ğ֟�B� ��0�N�T�f�x��� ������ү�>��� ,�J�P�b�t������� ��ο�:���(�F� L�^�pςϔϦϸ��� ��6� ��$�B�H�Z��l�~ߐߢ��6s5TO���/�#DO_CL�EAN�/�$6�NMw  �� a?��������g>DS�PDRYR=�p5H	I� `�@q�8�J�\� n���������������8��m8MAX�����17.X�-!*2|-!�"PLUGG0��*3�%PRC��B�^�b�'��Ox���
�SEGF� K���^�p�8J�\n���LAP �(�3���
// ./@/R/d/v/�/�/�/>�#TOTALPy	��#USENU�"; �8?�2s0RGDISPMMC� eo1C�@@@
�"4O�5 3_�STRING 1�	�+
�M�� S�*
�1_I�TEM1�6  n �-�?�?�?�?�?OO 'O9OKO]OoO�O�O�O�O�O�O�O�OI�/O SIGNA�L�5Tryout Mode�5�Inp?PSim�ulated�1�OutQ\OV�ERR� = 1�00�2In c�yclEU�1Prog Abor[S��1;TStatu�s�3	Heart�beat�7MH� Faul�W�SAler�Y_ oo$o�6oHoZolo~o�o�o �;�?�o�o );M_q� ��������8%�7��oWOR� �; o��oI�������͏ߏ ���'�9�K�]�o����������ɟ۟�PO�;�Q�����6� H�Z�l�~�������Ư د���� �2�D�V�ph�z����DEV� ��*���޿���&� 8�J�\�nπϒϤ϶π���������"�4�PALT�m[ч�5� �ߕߧ߹�������� �%�7�I�[�m���p�����I�GRI3  �;��s���'�9�K�]� o��������������� ��#5GYk��� R�m��}�� �%7I[m �������</�PREG_�H  �!/o/�/�/�/�/�/ �/�/�/?#?5?G?Y?�k?}?�?�?�?]�$�ARG_o�D ?�	����1��  	�$V	[
H]�
G�W+I�0SBN�_CONFIG S
�;IQHRCA�CII_SAVE  ThA_B�0�TCELLSET�UP �:%  OME_IO]�\%MOV_H8�@�O�OREP�_��:UTOBACK��ASMFRwA:\5+ _,5&�@'`�P5'dR�eC� q^ ,H5-�_�_�_�_�_*o]T���0oXojo |o�o�o�o5%Eo�o�o &8�o\n� ����S��� "�4�F��j�|�����p��ď֏��  PQ�SYSUIF.S�V ��R TL.�TMP XLED.GIF _$�6�8H�Z��ZqsAkA�0PINI^�5$�[E-SMESSA�Gw@���A�0��OD�E_D�@zFDV��Ox��ǟ-SPAUS'�� !��; ((O�2�1��Q�?� u�c���������������;�I����TSK  
�d__�0PUPDT����d���ԖXWZD_�ENB��WJ��ST�A���1���1WSM�_CFO@�5�]E�7�GRP 2�� 	BB� s A���9XISI@�UNT 2j��C� � 	z��� ��^ n�^� �� %�� �5*������ ���������0��T��W�i�MET� 2�u�PNߧ�J���^�S�CRD�1��P�EB��$�6�@H�Z�l�~�]_5*Q{I ���������(��� L���p�����������01�k��73QGRn���|�	UP_NA�@��;	3T_E�D��1�
 ��%-BCKED�T-���J��U /A�Uq4Rz5*,B�&o�Fs&  ��2�K�wʹ �E��	�-3�X5/|�/|/ ��k/�4�/$/ ?H/��/H?�/�/7?�/5�?�/�??���?O[?m?O�?6 LO�?�O�?�uO�O'O9O�O]O7_�Oe_ �O�A_�_�O_�_)_B8�_�1o���oxo�_�_go�_9�o o�oDo��oD`�o�o3�oCR S_���]��Ug���	 V NO_D�EL'GE_U�NUSE%IG�ALLOW 1z9	��(*��TEM*��	$SERV*¯�Ȁ�7REGх$�܎ȀNUM���	��PMUt���L�AY�Я�P�MPAL��J�CY'C10U�h�R�V���ULSUH�
�j���ӃL��ݔBO�XORI��CUR�_ʐ	�PMCNmVD�ʐ10~�>0�T4DLIȰß<�ˋ$MRߎ�&�&�ϲ����̯ޯ����y	 LAL_?OUT k���(WD_ABOR�o���m�ITR_�RTN�����m�NONSTOM ��� �շCE_RIA_�I������˰FF��U�c���o_LIM߂2` �  N��DNϯ�<��m�`���� ?Ϡϲ��ϯ��
����p��PARAMGP 1U��Ύ�O�a�s�>2�C>  CV���Ef��z�ߵߗЇ��U��Ж�Р�Ъ����Ԛ٢����������C���ǀ C�j���+���?�ɲ{HEC�ONFI��w�E�G_P�1U� 49������������E�KoPAUS�19� ,�uG�Y�C� }�g������������� ��1U?e��!�M��NFO 1�(�� ��=���� ������A�/����%q��w��Av��� D�a��q~D��Q�6������� ˰O����ǩ�COLLEWCT_�(��pEN`���\�I�NDEx(����!�1234567890��⁐�����H,��) '/L/�|&/8/�/�{j/ |/�/�/�/�/?�/�/ ?e?0?B?T?�?x?�? �?�?�?�?�?=OOO ,O�OPObOtO�O�O�:"� � ɶIO "��ǁ��O_a_s_�_WT-R�2#](�8Y1
�O�^P�$,]�Z���Y_MOR"�%� �9�Fe�Fi^o Lo�opo�o�kb�#�&-mB�?>�>��Ф�a�Kt�A�P�M(���a�- =�Oas�ϗ������^@
����` *c�P�DBO*���Ec?pmidbg�C�,��U�:��i)��p/���S�  ��фk�-�̏�������v����#������g�^�)� e��fM���w|���@ud1:˟����Z�DEF Y)o7S)ߑc�buf.txt���M� �p_L64FIX +�Q� ��˓�د��ɯ�� 2�D�#�h�z�Y����� ��Կ�ſ
��.�f��x�_E ,�  �l�~ϐϢϴ���p�+IM�C-�]��6���>���=L�-���MC&c.�SQdF�'�%d/5ݤ`�tձv��B!!� A*��B���B>�BZA�,BA���A�;�B���DB�"C���<C4�C�s�CC���D�2FB�n�E��E4���E���EC�2бy�bG��g1�\D��y**�~*�*�}��`U�xZ*�CÇЯ���BDw�4  E	�
��Ee�3Ec���Et� F��3E�ŚF��B� F���F��YfF�% G��� G	ڳH��3���  >�33 ;���aN�v  nf��q@�aG5Y���b�pA�a�t�<#�eDQ��7���F�RSMOFST '�f�GɫT1#`DZ�2!c���Q�*;�0��R�L�?���<��M��TESTR�0��FRz3S�Mx�C�A�z�D*e���| C�ЛB��C�pn9���*:d�b2�Iy4<2T_~�PROG ,k�%^�/%PNUSER  �1���KEY_TBL�  -e1]��(�	�
�� !�"#$%&'()�*+,-./�:�;<=>?@AB�C�GHIJKL�MNOPQRST�UVWXYZ[\�]^_`abcd�efghijkl�mnopqrst�uvwxyz{|�}~�������������������������������������������������������������������������������͓���������������������������������耇���������������������A� LCK#D#�STATi/0_A?UTO_DOG㺒��+INDT_ENB�/ �"��/�&�T2�/6STOP��/�"SXC� 2�5K�p8
SO�NY XC-56�Q{��p�@����	�( А{X5HR50�z�-tx?�>7�?�5ACff�:�O"O �? GOYO4O}O�OjO�O�O �O�O�O�O_1__U_�g_�\TRL� LE�TE6 �)T_�SCREEN }-jkcs���PU0MMENU� 16� < O\�o�u�_oIo�� &oLo�o\ono�o�o�o �o�o�o 9"o FX�|���� �#���Y�0�B�h� ��x���׏������ ���U�,�>���b�t� ������П	����?� �(�u�L�^������� ���ʯܯ)� ��8� q�H�Z���~���ݿ�� ƿ�%����[�2�D� ��h�zϠ��ϰ�����b��S_MANUAyL"?�QDBCO� �RIG�Ws)DBG�_ERRL� 7��[�����ߴ��� }O�NUMLI �I���dD
O�P�XWORK 18���&�8�J�\�n�DBTB_�Q S9<����K�,�DB_AWA�YW���GCP rD=����_AL �/��S�Y!0�UD H�]_q� 1:����0,R0�T�PA�~���_M� IS� ��@|� ��ONTIM�W��D����
�2#�MOTNEN�D'"�RECOR�D 1@� �<����G�O�N< ����z���G� �Nr'9K� ������� ��#/�G/�k/}/ �/�//�/4/�/X/? ?1?C?�/g?�/�?�/ �?�?�?�?T?	Ox?O �?QOcOuO�O�?�OO �O>O�O__)_�OM_p8_F_�_�NO�?�_ �_�_<_�_�_�_'o�N��(o_oqo�_�op�o�o�o�N���o �o9$2o�O ���&��\���5�G�Y����TO�LERENC��B�����L��O�C�SS_CNSTC�Y 2A~� h���Џޏ���� &�8�J�`�n������� ��ȟڟ����"����DEVICE 2B~� ��r��� ������ϯ�����)�����HNDGDw C~�Cz<�|��LS 2D\�;�����Ͽ�����=���PARAM� E/���?�)����SLAVE �F~�J�_CFG �G/�)�dM�C:\��L%04�d.CSV(��c�����A ��CH��n�n�)��=�[��)�-�Z�j�X�Wў�JPъ�C�_�CRC_OUT �H��<�+ϑ�S�GN I�����\�18-�MAR-25 0�8:33��)�05��16:01����� Ze��7-�)�)�*���o���Im��P�u�G�=��VERS�ION ���V3.5.20���EFLOGIC� 1J% 	���* ������PROG_ENB�����ULS�� �,P��_ACCL{IM�������7�WRSTJN`����)��MO��
��x�INIT cK%
��) v�wOPTp� ?	�����
 	R5�75)���74��6J��7��5��1�2���6����TO�  ��@���V.��DEXd�d��x���PATH ����A\����IAG_GRPw 2PI�|O��	 E7� E�?h D�� C�� C ��B���C��n�k�����C���Cm�B�N��BzoOB�)��Bk��f383 6789012345����B�  A���A���A��A�O�A���A{+A�s�Aj�RAbJAY%, x�@���p��G!���A�����BA4h���x�
"�����"�Q�A����A���A߈��A�� ���hAx~�Ao��7Af9X��?$>��mF/X/��h�����("_�AY��;AS�TAM��^AGdZA@��A:bA3�%A+�-A$���)�/�/��?�*�@�;d�6����@{�@u�-�@o�@i�7�@cC�@\�j�@V{N?\0�5�?b?t?�??@_���@Z^5@T���@O�@IG��@C33@<��@6�+@/<@(�`J?\?�?�?O��8s� nE�@h��@b�!@\��0Vff@Pt@I�hs@B��@;�bOtO�O�O�O�' 6]^_p_N_�_�_0_z_ �_�_�_�_$o�_�_
o lo~o\o�o�o>o�o�� C"�!30�2KA�@^�>8Q�r��R�?�  *u^7��ŬFr'Ŭ5A�FRu^@�p��nv�@@�pppE�@�[ Ah���uC=�+<��
=T���=�O�=��=�<����<�p�q�xG�� �?� �C��  <(�US�� 4jr�D@���Y�"�A@w�?f �oX��mf�������� ��ԏn��
��.�@���i?#�
b���\>�pn�^��G���G�^x���R����^8�ۑ�5����CnB��L]_u��&�
P;�'f�d��aQ�{���dD�  D�  C΍��̯ޯ 8����@V�ǯD�ïh�������3*Da��q�D�Q�7�f/´�S�Կ w������.��Rρ��!�'��t�>�6��=ݠ?�8xA���m�Yϧ� CT_CONFIG Q-y��#�c�p��� STBF_TTSd�
����C�tV����MAU^�����MSW_CF���R-  ]z��O�CVIEW�SY�i�����߽��� �����G��.�@�R� d�v��������� �����*�<�N�`�r� ����%��������� ��8J\n�� !�����" �FXj|��/�����//j�R%CR�T�e&�!�,. V/�/z/�/�/�/�/�/��SBL_FAULT UI*n�1GPMSK��$7���TDIAG V���e���1�UD�1: 6789012345�2��?�P�Ͻ?�?�?�?OO )O;OMO_OqO�O�O�Op�O�O�O�x �>��;�
�?%_��TRECPZ?l:
z4l_?� �?�_�_�_�_�_�_o o0oBoTofoxo�o�o��o�o�o�O_/_U�MP_OPTIO1N�>*qTRR���:!9KuPME��>�Y_TEMP  È�3B���p�A�p�tUNI�7��şqF�YN_B�RK WY�)8E�MGDI_STA`�u&��q ��pNC�s;1XY� ��o7�*�~y���d ���� ��Ǐُ����!�3� E�W�i�{�������ß ՟����Xu"�4�F� X����f�������¯ ԯ���
��.�@�R� d�v���������п� �����%�7�I�[�u� ϑϣϵ��������� �!�3�E�W�i�{ߍ� �߱����������� /�A�S�m�w���� ����������+�=� O�a�s����������� �������'9Ke� [������� �#5GYk} ������ /1/C/�oy/�/�/ �/�/�/�/�/	??-? ??Q?c?u?�?�?�?�? �?�?�/O)O;OMO g/qO�O�O�O�O�O�O �O__%_7_I_[_m_ _�_�_�_�_�_�_O o!o3oEo_Oio{o�o �o�o�o�o�o�o /ASew��� ����_��+�=� WoI�s���������͏ ߏ���'�9�K�]� o���������ɟ۟� ��#�5�O�a�k�}� ������ůׯ���� �1�C�U�g�y����� ����ӿ���	��-� ?�Y�c�uχϙϫϽ� ��������)�;�M� _�q߃ߕߧ߹���E� ����%�7�Q�[�m� ������������ �!�3�E�W�i�{��� ������������ /I�Sew��� ����+= Oas����� ���//'/A7/]/ o/�/�/�/�/�/�/�/ �/?#?5?G?Y?k?}? �?�?�?�?���?O O�?K/UOgOyO�O�O �O�O�O�O�O	__-_ ?_Q_c_u_�_�_�_�_ �?�?�_oo)oCOMo _oqo�o�o�o�o�o�o �o%7I[m �����_�� �!�;oE�W�i�{��� ����ÏՏ����� /�A�S�e�w������� ��������3�%� O�a�s���������ͯ ߯���'�9�K�]� o���������џÿ� ���+�=�G�Y�k�}� �ϡϳ���������� �1�C�U�g�yߋߝ� ��ɿۿ����	��5� ?�Q�c�u����� ��������)�;�M� _�q�������!����� ��-�7I[m ������� !3EWi{� �������/% //A/S/e/w/�/�/�/ �/�/�/�/??+?=? O?a?s?�?�?�?��? �?�?O/O9OKO]O oO�O�O�O�O�O�O�O �O_#_5_G_Y_k_}_ �_�_�?�?�_�_�_�_ 'O1oCoUogoyo�o�o �o�o�o�o�o	- ?Qcu���_�_ ����o)�;�M� _�q���������ˏݏ ���%�7�I�[�m� ������ǟٟ��� �!�3�E�W�i�{��� ����ïկ����� /�A�S�e�w������� ��ѿ�����+�=� O�a�sυϗϩϻ��� ������'�9�K�]� o߁ߓ߭��������� ��#�5�G�Y�k�}� ������������� �1�C�U�g�y����� �����������- ?Qcu���� ���);M _q�������� �	/%/7/I/[/m/ /�/�/�/�/�/�/�/ ?!?3?E?W?i?{?�? ��?�?�?�?/OO /OAOSOeOwO�O�O�O �O�O�O�O__+_=_ O_a_s_�_�?�_�_�_ �_�?�_o'o9oKo]o oo�o�o�o�o�o�o�o �o#5GYk}��_ �$ENETMODE 1Y�U��  �P�P�U��{��pRROR_PR_OG %�z%�V��&��uTABLE  �{oe�w�����w�rSEV_N�UM �r  ���q���q_A�UTO_ENB � �u�s�t_NON΁ Z�{�q��_  *����%����Ā+�*�8<�N��HIS���Q��p�_ALM 1][�{ ��T��P+O�˟ݟ����%�S�_����  ��{��rj��pT�CP_VER �!�z!�5�$EX�TLOG_REQ�k��ቼ�SIZ\ů��STK�������TOL  ��QDzs��A= ��_BWDJ���؆K�ԧ_DI9� \�U��t�Q<�rU�STEPa�s�|�p��OP_DO���qFACTORY�_TUNk�d̹D�R_GRP 1]�yށd 	e�#��p��x����� �n��So �k� ���W��i� z�dϝψ��Ϭ����π	����?�*�c�N�@�p�@��?���@%:�j�
 F�5U����j��xd����E7�� E?p D�٠��L�D�%�� � C���K�B� } ;�  A@E�^o�@UUUc�U���K��w>�]�>�y����ѻ� E��F@ �ѿ�{�L����M��J�k�K�v�H�,�Hk�{��?�  �Q�9t�Qv+�8���6�h�%7�{�]�� p2J��1����/ �j� g�,�FEATURE ^�U�K��qHa�ndlingTo�ol �� rod�uChine�se Dicti�onary��LO�AD4D S�t��ard��  �NDIFAn�alog I/O~��  d - ���gle Shif�t��F OR��u�to Softw�are Upda�te   J70� matic B�ackup��ar�t Hgroun?d Edit����708\��ame�ra��F��D p�r��nrRndIymM��PCVL���ommon ca�lib UI /q.pc�nf� Monitor��owset�tr��?Reliab	 ���jp Data Acquis������ Diagn�osD����� D�ocument �Viewe����
PC ual �Check Sa�fety� ac�t.Enhanced UsG�Frw ��\weq�pxt. DIO� � fi+ t\�j7�endxEkrr� L*  � ��{s  ��r��� :���T "�� FCTN Me�nu`v���t }I�TP In��fac%  48�\� G_ p Ma�sk ExctgԄ� o��T Pr�oxy SvH � 5p��igh-wSpexSki� " #1��#��mmunicC o�ns�apd�!u�r �����"c�onnect 2�Pdin� ncr� stru�� �I KAREL �Cmd. LE u�aG"t\ia�%R�un-Ti�En�v��"K�el u+G sE S/W��Licen8��[GER  ��Book(Sys�tem)�� R5�� MACROs,�x"/Off� �P�a� MH�- �: 7\ac�1MR� ��)��MechStKopV!t�  ��0i���Mix�x��E ��
� �0o}d
 witch��GLoa� �4.�6� k G�1�3Op�tmUHM GGW fiIlG� HF��g�'� pmfO Mul�ti-T= i�4p�a�PCM fu1n�'{3M"Po[��D QV�HReg�it0r�   mp]o� Pri@F�K� _fcs W g Num Sel�5���� DS� AdjAu� ���`W
 4 =S|XtatuQ/�bUC�� RDM Robot���scove�� c;ctO Rem�0��n���SServ�H10@#CTXP?SNPX b<2��� "K9$`Lisbr���564@eb�� �4H`ZUSoY0=t ssag�E��~� "�1�VVLO��b/I- pc}
�`MILIB�m�ch1o Fir�m+�8� �b"Ac�c` hXcTPTX�;��� s Teln��0�m}B��5��4T�orqu
 imu�la�}�Tou�7@Pa51��m�T�_ �QC&V ev.� ocleU�SB poU � i�P�a@WdUSR� EVxP+Un?exceptx�P��D{D{f}VC�r�"�"�2�sVD��jx�cV�Hk uifo�V�SP CSUI��k��XC�6X`?Web Pl�V���9pjăa�+64.f��^ r>�T�vΛ
J57À�vGr�id�Qplay 76 (��`L&KiR;�.��K�\0�ARC; 4 120�i��L#Ascii�V!eRDAG�d��Up�lE@��� �@Col�lW�Gu�� of4^QޝPI   1�s� ��t�0t8FK����Cy�p  2*Por�ie  ld�aF�RL�1am͉ R�INT��MI D�evO0 (&ax2 �,�0�%(}t\rb��A/��Passwo��:O" {ze�s�
! 064MB DRAM�
�qG`��FRO�� �RBW��rciPv3is�]�BW� .��Welds cia�l�4 "P��el�l���mrw�s�hg�s���cXE aSwm��( p�v �Q���ty	 sPR-�8��2�t!1m@.�bo+�D�P���D� 2b a���r�Dr��Pb� q ged�� rT1� e8sOL��Sup�r�AR� ! � OPT �"W�  ���; cro�V ���SHe[��;`L�Qfq�X�ueOst E�$`S���e�tex{DSAp$![��P�`P@ �4YF�VirtxW�S��  ���stdpn�x�u�io SWIMEoST f� F0����&�� аߕ��51 J����(F9r�ߕ�II)�ߓ�on��!���M!=��RY���f>�t���mfV��լ���Ҍr�� ��?���&P�3����Ҭb9���eie.T���n\p���\R���ҭ`A��2�p�����!
!����O<����7 J5�����5�ӝ1Q��\a�r7���XPR���k "��}��b���r�`P���lnko�0i���0��RMJ�Ո��;���M�����Hs54���j883�]DER�N��Ffh�M/el���չ1d/������d0�/ ��|B�/�( �/��<���/��p��?��.f9d�/��ASTC?���616�/��g HaS|?z��as��@����M��?��0�?c�r W$O��!`���%rzP]O��t\awxOV4�`�O�$�a�O �ҵ��O����O��.�EN _�D�`<_��i�te_?��v �t_�� aO=%IF�{?�Ԉ`���) "�s_�Epa�O-�>n1�!Ot.vTo5!��_��F���o^83!7�o*QogW-���o��/5-X@�PDT`4B��Q��ze�O2Hf4�_\79���MN������f�t!ro9?6�x�i0��ԇJ59L��%����A`k��P����_p�o�Fp_-o�@�?�(�f1'?�pm_ d��O��ٟ�O.�3pe����m\�A���/_����2.p�͆cW_�֮͠c�8a/\ R8���(Las$���O_0���0x���bo��<� ���e�̿"% ���8K��/?�sif<Ϟd��?�NT+���Se ����//�C/��̕��'37��iUf\�����$SG��Ԁ63q��RDYLS߱��oI�omw��_#�p�s0�����hVmLj��93����E�o@gW�P��ch\?�I��ퟓ� �o����'rvi7�]S�/��8����V(st,��F���@�tl�u&5�/����T
�hWi��ݶSe��6O��csr��	��! b��y8P`�dr׏��o3PRI���a��O�/	X/��s�pr�ߕ����Li<?/��3 H6x/�d�94'��63�q54s H�/v653�/&r4 H���&0�/�'`��� X?v72��Ie?�g13;?��7$�/58r?�'6�/��3Lo�_��t �ͅ`A�ϐOc�m�osK� !����O����,�O9�8�O�OS�ualP_���8�?a_�^��<̤_��wr+��j8�3�?!�_]���ND$SO-�f7O=�!�Y�3ad�O9kl�o�s_#1�o��ip#�-E9t�op�RIN,��3/I���VA�=�SE_��0
S����Z 0+ͅcmg�Z�� 4@�"�ut[/�of��`��M�r����@����5�96O_��4Џ��U���#o(� I�c5%rA_����e`���G��������c��AL9"���lg33_U̻oy� -<�t
௟	e�@t���RTU����h�z�xo��vao;��'O�52 @����4��'�Yu\��F vOA���4I`FĿ&
d -�ݕE���c (o�[�"E3�yo��Wel_��������WMG�Ϣ3a8P@�Ϣ3wmg[����߂�- ���On�345�?�fCMk�IO��  �ߪ�������1���2�g�y� R��;�Co���4(S�`�⯔�Ġ��33IF���� !(�z�f0at��NT��q���R8��i5�P�g82\��� O ��W?��˿ݿ￘��7��4SiZ/<��=��K�!�cl�i5\s�w/�S�AD���C�Vt�Dt.�Q�m�t�_�e���V�-V0�  /6��Nlo��1"��\�O�/C �/�4 �/�i�e/�/L1_��62˟��o�/��eJ7��erv��?�) "�?�svh�?
o�N� �?�s.p[�tvhmoO�U749LOR`r���OutlO?�t\�?��j�_�//�/�h_ mpc��y�9	\KO�j�_�/�_f�uXP�/D�H8gOL}�oOnn�O�%N�� �u�'o���n]`���NoRCM�o�un�_ ��$./_#���m  Hw552�abe�q�38BSR78�p�q�r0��lib�J614�c�ATUP�@rm�c�p545zPsg�t�r6�VC�AM�3CRI��p\rc�pCUI�F�  �q2�ptd�.f�NREN r�co�p631  �- Pr�pSCH�V� DiDO�CV>aIFL�CSUUJ18�0�p1}��EIOC  Z��4�p54�pR�`�4�9�pgm�SET�f�Sta�q�qla�y,�p7�q�0�MASK�SoPRXYZaap��7f�C�pHOCO�C��3.3�r�p\c�΂51�p��qap�p.�q39f�j5�0�q�ust3�L�CH��A`
O�PLG�1"�E�� �"L3�MHCR _ 08 (ĀS@�7Reg��CS�p�1�H��p��q5�p08�\�pMDSW  7URGw�MD���s�OP��\!�MPR�ra�4�Հ!�o�f���p! p��PCM��H��R0БPa�th���p@aH�ՀR�m����pTP���Հ8[16�50�pg���āS��ol,�9Ղ:�FRD�p(Q�p�MCN��cc�H�93�pLNP��S�NBA@�rSHL�B��֑SMx�lr�n?�63�p��q2��pL�HTC�pX�TMILVs�r�T���PAu�Y�sȡTX�>aEN��ELU�tEh��0�@`�8�q`HѰr9��`ρ95�p� �Հ7��UEV^��adin(�C��ܵ��pUFRI�ee�O�VCC�pt�VC�OY���VIP��s�pd�[�I^�p�Xv͡tsπWEB�p���?�HTT�p L�2�R62�pCoo�?�CG��d�I�Gt�
PRI��P�GSN ng�IR�C��ne ��H8m4�prd6�R7���@�R��L�53�p\�lcl�q8�pD"� #4�6M� ��592�8�R659��:|�5�r dK�6��p��4�49�YpS��pp5�̰T©qG ML��06�pg, ��F�{���ð��pJ64�3�pWS�p��CL�I�zdҡV��pGD����u�$������h�TY��<q�TO�pg���q6�-@��sR5 ��ORSY��3��68�pģOL�p�sguK�OPI�ɰݠ�pS5�R�RL�P�y��S�2!�E�TS1���43 m!��CP-�ryB��VRu�onF�IP�N�� Lo��Ge;ne~�(SytE�a��I�0�՘��p��ytt\sg��g ="�ր6q��L�yt\str�ոA��<�A��hk_t���yt����es�լr��{j7��mon.��(�A��d@6��s-@����yt46\�`Q����qh3��zDlli�4�F�lc�`�$rt{���¥���yt��w�x�U�Ӑh8��nde��AxV絰�����N��ͰH��epCen���yt�T�ՌĢ��ob3攢��hS89����p��Pv�sed����4 J7/R805��0l���:�`"t644������ II���r�p����"S��5л%���594G�tomt���!�R J�ؖ� ��Se3�ar3�E�t32�%�QsysG�F ���������etr��ur1nk����20�xc78���'�rn6������\jtET��
jo��ta.C����gr������`� ���<���ge�.��017��2�ytL�yt75b���Lj(t���7 "P��T`dc��) ���	����r��1%a�t�@O���p��daW(?�4tv/ 4oh��c8}���s?yR�?��=logm�?�;ild�?1<d�?N�@ ���0@O�M���p1|O�;x@���ytV�B�1���O_�	8�7aicC 2�9���C��7��6o�E �� `�E?kedg?y=wm�`ORhl$_�2G&�he>�m_��7�5�l�O 24O Oaw�4OJmdh\o�;dhq2���osqz�o�kl���o�o��:��+�F�et�'-�6J�8"WQ��1 (F����pDa�0��f�r{F� �� �f22�.f�FusS�pkYg�M!INgD�x���,��u��o�{Ώ�522�xsiR=C�n VM��^��992�W� ��J9�b�st�'T��Oo 92\�6CMR/@d#Z��O;��ݎv'�D��tmF����f8��vat��t+9�>e��6ft"/��zC_v(��ɟ?�4o "��,���կK����cvsw�8��Dni�o��lb��蟮������W�\���vsmTڴaz�"����ο��of���1ow�(ώ�slw���f���e�w�����*ԣvr�ys�+N3Ge�N���Y25:�oa]d��(Na�NJ�?��nd�� "N�wV  �@��s<���rrd�6`��le&���C�bU�4;��Ok7\���8���rk&,��gl���P��g�Gt��i�l������  � P2^���38��r �����0��J61�4�ATUP�j���545����6~F�VCAM��_CRI!7� N, UIFB���2���ans��CNRE��'��631��RI��SCH�u65�DOCVN�ns�� CSU�T|���0���HAEIOC�% "��54��R�6965\� ESET�W������7 Cu� MA�SK�t 1/PRXYUJ N �7�ל�OCO�o]m�513r�,,������� ��98\t�����]�[39�v!���oftw�LCH!g�OPkLG:�950a�i�P]P��e f�,S�r��CS����g_lo���5� �pDS�W6�r70<!Pl DKOPP4�;PRQS01� n �Ad����X#PC%MAa ��0�%���vdv; �A
TX��0��1ADIG� ��!H ,S�r72�3��9AU�+ FRyD!h#RMCNr	�H93��R2SN�BA"�C+ SHLB�	SMp5�n �m�J52�HTyC���TMIL6ԣSe���PO�0P�A�86*TPT�X�VR�0ELA4oGol,��� P��8��\sv���qoSRVT��95Qv$95A\et� GUEV�@a\AC!,]�[AFR!r���C!ol.�VCqO��P��VIP�4ie�� I�t34[�SX���WE)B���@(�1T��,��l2tQ, G�Eg[\tkIG�E#@`�PPGS"�PRC��4"TAN��84l��#R7�taQ�R�(
R53�t�RJ68��R6�6a52a- �E��R65qr Im�5a��l��w573R64q���q5`M�RQ�C�D06��,0g�  �R40�AAkWS!f9LIq%�ni�@�P�SCM]S�597[M%o76 J\0TY�4�L�, TO��9 (vk76�fer@sR5PCORS�w\snKR68��CSN� ��Eq��=I1Tcsn.\0� 6��cL�EX�[1�f��� TS1Th#� ��P� �0a �,0VRh��,QN�4Ca
AGeneH抳�y�MG" �y���yg�_cc�y"�xcm�g_�y��yvth�yR�x3(�,�>�P��b��z1��z! cv�yon T�yh"�xhr�x�b݉1�`]�iA��y CV�yCP  �z��x��xt���	q��ypse������r;57� In���w�x͉576��(p�+�)� ����L� "yAl��w6\ab����j8<�B��h ���PR<�J8�zPcxC;�8�J�ps��9P��x96\{�(P��y�����A�x9 � �-��iv{�R DmM<�H7�zH6�{66�3�1�x�[�tor�������y�m�!��sZ�]�92����nalۺ�Й)�޸stK��}s3tr��ypsk���=�\p����xj932|�C��}�)��x8R�x2}�����.�|�޸_w���}hk�_k�FH���9!�xk5e*�n�95
����yhe�z��<�,�f�l.��H�eGt_w�y�"M�c� �� �zbak�H�Z�gent��h�\m���s���� ��d�� ���Y�;�(�Z�@�z
9Pf�yv�@��.��� ��� l�n�( l��gd��=
i��! xZ���+�00iB\��H[�H���� -�h�[�C" #��822��2�@}�OR��� ���iB/̿N@�"F���f��h@+�t=���tk� OR��ƈ�83�i1�t �˚�~nc+��fc䫚��5���835 �z����i�;�5:�B6�ri��ER���bv݉ (ˊng,�@�,4�*RȭY��k=�mo�`]/��p��+��ptp�z(�5\pk�=O?����0[� ���0�/�/ ?S�i�k߽�ij��
��?�+��db��� s5E0l�a��x���S�[�d G�yϋ�ce���0K�50�K1^�y�6q�Je��RDE��yqInt��
 Pa��(�9\9g{�H�919[�pܻ\:� Vi��to�ol<?ވ	�J[�ucppK/=_��vk{� �K[��Z��Z��O�O��O�8�OK�H��?�G_srj;*h�ndr{�NH]end��Ir:�b(�3��o~H73;���/�&7;*��{X��j�|���"�4�  �am_xO�veH�ʘ���vI���o�?�|�xj{��� �T�z{�] R5;�J9�;989ﭹ���_��p�m
�
�`��:��e�kR R�}++�R7�J L:;) !"���Kz�/p+zx��d	�-�|�	�63=3�06 S�I~R6�st�z��:�wLND��IF K�s45��-con{
qC9�i�*ar �jxyp�	�ds "�����ENl�y��sl��l�gr��e-�
���856��`�zr�piZx=H�4� l�^�wj�! r6˛vv�:nn�}�RC:| �� J9��Z����867�1E3J;6��8 �JT�`��I(iR��R|"�ٟc  �STD��.p�LANG&�����r��ti����P��q���)0-�� E��kgS
��y` ��5����R730��(���8 (i��ErreP��,�`��PC��<x���rvge������8���ge��a<舰��	�.��isi=o��ckin�� ��R�(���pGi@� �����؁��j	���PFK"��XA��9\@��BP4��!x��d��aabbPbbb�����P��P��(1��SP�Р��FS J��J91.��6859!	�֠�02*4<62�7���Y��,`����X���s\��GFSO����scex��/�vr��`���&���RG(WR68'64��p���#8	G (� CCR��I���;cc�� "CkH����9�\RBT�}rgOPTN�4�4�2�4�?�?O^"Ocrg.8EF���8E��
8Ed�D{PN��ion �E�nd.�Exa�FI�NT�E��7�E� n"�Ea�@�E�0"�EHQހEhd\m�FHDx�F��D\erh�F���O�Ai�E��s@BT�!Uire�Eh�Dt�Drh�GdCfU��ted ��-�n� An�U��-�9p9 �Ut2-�8-�0E-��a�U�`t f�1-��2-ĥ m�U�a�U葬U�-`s�U�ѬUpB-�1��-Ā6q�U wR88�U851_fy4�`�Utiar�U�-�it� -�l"-ďMR S�f`�fTcXP�U��epm�f�" #1�f! T�fy��fm�g��e�P��U 2�U 70�Uo�njg-ĭ@_f J�7�Vipp�fon,��U���X�v4-�j7�9�fc��e]h98xjg�"-�\chp�W�EN�vd@Pb{St�o'�� E f�@�VgF0�el�gxѬU���j8svY��f�-�6�uharel�UKA�Ro�Comc�u�R�ĆL*wp\ �V
t+vY�u�fp\e�V�AN"���k�gpcp_f1a!I�[�f�4y�wf
! Gf ;Co�uarwf��FІ84_f5 H�fH84�v63 �H�fH7�v779�_f24��7rw69V*�65�f1�g8p�v�V75�VIC �fw AP7v893�`��R0-��B�eck���Hs�
E����#fMNS+v���VՐ�V�P_f-]�_�Q�V8X�\���tch믅��U3\pSfWT"p_fdBe��Zhin_�� �03jgoXЬU(7ROB�wOG���A�Ue�A�^�HR�Px`flRuuyQuug_Sfz̉3uh523.�U{le*writy ��6�2�6�5sv554f�4І40����H60�v0�h�[�08��+�=�O�a�b��8< ���68v�`��s�75^0��A�rw7��h����וл��3�v3Y� &�U �େ2f���� 29#f�p����\ib<f��;sbs8�w��o scbP1o�Cja��Ly2%� -k�E"�74�V9 wf� (W_�	`��XPLF���wvF�E�X�φ�`we�Vp��a\cwvTf͸�z50+�G"WV����֤u���2�Y �� ��nte�g�����f04 (��gx��D����BP	Xk���I/��`o�!d�@��G��pv �kϥ�ib�hp 
om �wfE�A�f��&Hfdn���z8Z�0f��ؿ�ra�W�_��oi �<�al�VV�Ax�V�2�� 996#fVCA��,�vast#/�q� ��"��dp/fyn:�f�i���58����D��odif��.e8�DP��q (d��o "���o��Rg�d98Ԑ'G��strS����OAW���wR73��v16"� Rf�7�9�2���iTra���c�h�/�wv"�TP+v̀��tpe��c�wor���+R�C�59�8�� S�5+�809�?��C��f�"z\mߦ����RE��$sFL&0�pcz��6�verv�gng�_��746�_��S�_� Ch�?�� {�����<t�h��0�897i3��g����:�f!Ě��Īx���� T��w& ���rk����`s��H�VAGǧset�99�b����$FEAT_A�DD ?	�����q�p��	 x������*� <�N�`�r��������� ̏ޏ����&�8�J� \�n���������ȟڟ ����"�4�F�X�j� |�������į֯��� ��0�B�T�f�x��� ������ҿ����� ,�>�P�b�tφϘϪ� ����������(�:� L�^�p߂ߔߦ߸��� ���� ��$�6�H�Z� l�~���������� ��� �2�D�V�h�z� ��������������
 .@Rdv�� �����* <N`r���� ���//&/8/J/ \/n/�/�/�/�/�/�/ �/�/?"?4?F?X?j?�|?�?�?�tDEMO� ^�y   x�=�?�?OO %OROIO[O�OO�O�O �O�O�O�O__!_N_ E_W_�_{_�_�_�_�_ �_�_oooJoAoSo �owo�o�o�o�o�o�o F=O|s �������� �B�9�K�x�o����� ��ҏɏۏ����>� 5�G�t�k�}�����Ο şן����:�1�C� p�g�y�����ʯ��ӯ  ���	�6�-�?�l�c� u�����ƿ��Ͽ��� �2�)�;�h�_�qϋ� ���Ϲ��������.� %�7�d�[�m߇ߑ߾� ����������*�!�3� `�W�i������� ������&��/�\�S� e�������������� ��"+XOa{ ������� 'TK]w�� �����//#/ P/G/Y/s/}/�/�/�/ �/�/�/???L?C? U?o?y?�?�?�?�?�? �?O	OOHO?OQOkO uO�O�O�O�O�O�O_ __D_;_M_g_q_�_ �_�_�_�_�_
ooo @o7oIocomo�o�o�o �o�o�o�o<3 E_i����� ����8�/�A�[� e�������ȏ��я�� ���4�+�=�W�a��� ����ğ��͟���� 0�'�9�S�]������� ����ɯ�����,�#� 5�O�Y���}������� ſ����(��1�K� Uς�yϋϸϯ����� ����$��-�G�Q�~� u߇ߴ߽߫�������  ��)�C�M�z�q�� ������������ %�?�I�v�m������ ��������!; Eri{���� ��7An ew������ ///3/=/j/a/s/ �/�/�/�/�/�/?? ?/?9?f?]?o?�?�? �?�?�?�?O�?O+O 5ObOYOkO�O�O�O�O �O�O_�O_'_1_^_ U_g_�_�_�_�_�_�_  o�_	o#o-oZoQoco �o�o�o�o�o�o�o�o )VM_�� �������� %�R�I�[�������� ��Ǐ�����!�N� E�W���{�������ß ������J�A�S� ��w����������� ����F�=�O�|�s� ���������߿�� �B�9�K�x�oρϮ� �Ϸ���������>� 5�G�t�k�}ߪߡ߳� ��������:�1�C� p�g�y�������� ����	�6�-�?�l�c� u��������������� 2);h_q� ������. %7d[m��� �����*/!/3/ `/W/i/�/�/�/�/�/ �/�/�/&??/?\?S? e?�?�?�?�?�?�?�? �?"OO+OXOOOaO�O �O�O�O�O�O�O�O_ _'_T_K_]_�_�_�_ �_�_�_�_�_oo#o PoGoYo�o}o�o�o�o �o�o�oLC U�y����� ��	��H�?�Q�~� u���������׏�� ��D�;�M�z�q��� ������ӟݟ
��� @�7�I�v�m������ ��ϯٯ����<�3��E�r�i�{�����˽  ¸��� �)�;�M�_�qσϕ� �Ϲ���������%� 7�I�[�m�ߑߣߵ� ���������!�3�E� W�i�{�������� ������/�A�S�e� w��������������� +=Oas� ������ '9K]o��� �����/#/5/ G/Y/k/}/�/�/�/�/ �/�/�/??1?C?U? g?y?�?�?�?�?�?�? �?	OO-O?OQOcOuO �O�O�O�O�O�O�O_ _)_;_M___q_�_�_ �_�_�_�_�_oo%o 7oIo[omoo�o�o�o �o�o�o�o!3E Wi{����� ����/�A�S�e� w���������я��� ��+�=�O�a�s��� ������͟ߟ��� '�9�K�]�o������� ��ɯۯ����#�5� G�Y�k�}�������ſ ׿�����1�C�U� g�yϋϝϯ������� ��	��-�?�Q�c�u� �ߙ߽߫�������� �)�;�M�_�q��� �����������%� 7�I�[�m�������� ��������!3E Wi{����� ��/ASe w������� //+/=/O/a/s/�/ �/�/�/�/�/�/?? '?9?K?]?o?�?�?�?|�?�9  �8 �1�?�?	OO-O?OQO cOuO�O�O�O�O�O�O �O__)_;_M___q_ �_�_�_�_�_�_�_o o%o7oIo[omoo�o �o�o�o�o�o�o! 3EWi{��� ������/�A� S�e�w���������я �����+�=�O�a� s���������͟ߟ� ��'�9�K�]�o��� ������ɯۯ���� #�5�G�Y�k�}����� ��ſ׿�����1� C�U�g�yϋϝϯ��� ������	��-�?�Q� c�u߇ߙ߽߫����� ����)�;�M�_�q� ������������ �%�7�I�[�m���� ������������! 3EWi{��� ����/A Sew����� ��//+/=/O/a/ s/�/�/�/�/�/�/�/ ??'?9?K?]?o?�? �?�?�?�?�?�?�?O #O5OGOYOkO}O�O�O �O�O�O�O�O__1_ C_U_g_y_�_�_�_�_ �_�_�_	oo-o?oQo couo�o�o�o�o�o�o �o);M_q �������� �%�7�I�[�m���� ����Ǐُ����!� 3�E�W�i�{������� ß՟�����/�A� S�e�w���������ѯ �����+�=�O�a� s���������Ϳ߿� ��'�9�K�]�oρ� �ϥϷ���������� #�5�G�Y�k�}ߏߡ� ������������1� C�U�g�y������ ������	��-�?�Q� c�u������������� ��);M_q ������� %7I[m� ������/!/ 3/E/W/i/{/�/�/�/ �/�/�/�/??/?A? S?e?w?�?�?�?�?�1�0�8�?�?OO 1OCOUOgOyO�O�O�O �O�O�O�O	__-_?_ Q_c_u_�_�_�_�_�_ �_�_oo)o;oMo_o qo�o�o�o�o�o�o�o %7I[m �������� !�3�E�W�i�{����� ��ÏՏ�����/� A�S�e�w��������� џ�����+�=�O� a�s���������ͯ߯ ���'�9�K�]�o� ��������ɿۿ��� �#�5�G�Y�k�}Ϗ� �ϳ����������� 1�C�U�g�yߋߝ߯� ��������	��-�?� Q�c�u������� ������)�;�M�_� q��������������� %7I[m ������� !3EWi{�� �����//// A/S/e/w/�/�/�/�/ �/�/�/??+?=?O? a?s?�?�?�?�?�?�? �?OO'O9OKO]OoO �O�O�O�O�O�O�O�O _#_5_G_Y_k_}_�_ �_�_�_�_�_�_oo 1oCoUogoyo�o�o�o �o�o�o�o	-? Qcu����� ����)�;�M�_� q���������ˏݏ� ��%�7�I�[�m�� ������ǟٟ���� !�3�E�W�i�{����� ��ïկ�����/� A�S�e�w����������ѹ�$FEAT_�DEMOIN  �ִ���ΰ��INDEX������ILECO�MP _���7���-��SETUP2 �`7�A�� � N l�*�_AP2BCK 1a7�?  �)Ҹ��"��%����ΰ:��� ��Ե��*߹�N���[� ��ߨ�7�����m�� ��&�8���\��߀�� !��E���i������ 4���X�j������� ��S���w���B ��f��s�+�O ����>P� t��9�]� ��(/�L/�p/�/ /�/5/�/�/k/ ?�/ $?6?�/Z?�/~??�? �?C?�?g?�?O�?2O �?VOhO�?�OO�O�O QO�OuO
_�O_@_�O d_�O�_�_)_�_M_�_ �_�_o�_<oNo�_ro�o�o%o�o�oF�z�P�~� 2��*.cVR�o�`* �F�cLpZepPC�x��`FR6:D��~\��{T� �'��u�Q����w�Yf*.F
���a	�s��Ռd�����STM �"�-��p��Y��`iPe�ndant Pa'nelY���HO����?���[�����GIF�6�A�"�ߟ񟆯��JPG����A���0c�u�
��zJS�=��`У+��%
J�avaScripti���CSZ���@����k� %Cas�cading S�tyle She�ets�_`
AR�GNAME.DT�lD�\0��P��`�q��`�DISP*g�J�D����σ�����ϡ�	PANE3L1��O�%D�8�x�k�}�+�2m���b� ��~ߐ�%�0�3��W�@b�E����0�4u���b�����-�(�T�PEINS.XML4���:\H����Custom T?oolbar�����PASSWORD���}nFRS:\����� %Pas�sword ConfigXoV�� O��o�?��u 
�.@�d�� )�M�q�/ �</�`/r//�/%/ �/�/[/�//?�/�/ J?�/n?�/g?�?3?�? W?�?�?�?"O�?FOXO �?|OO�O/OAO�OeO �O�O�O0_�OT_�Ox_ �__�_=_�_�_s_o �_,o�_�_bo�_�oo o�oKo�ooo�o :�o^p�o�#� GY�}���H� �l������1�ƏU� ����� ���D�ӏ� z�	���-���ԟc��� ���.���R��v��� ���;�Я_�q���� *���#�`�﯄���� ��I�޿m��ϣ�8� ǿ\������!϶�E� ����{�ߟ�4�F��� j��ώߠ�/���S��� w߉���B���;�x� ��+�����a���� �,���P���t��� ��9���]�����( ��L^������� �$FILE_�DGBCK 1a���� ��� ( �)�
SUMMARY�.DG�hMD�:�0t Di�ag Summa�ry1>

CONSLOG&	t��CConso?le log�=	TPACCN��/%�4/?TP� Account�in�>
FR6�:IPKDMP.'ZIPh/l
�/�/�@P Except�ion�/n+ME?MCHECK*/��@?�Memory DataA?��LN�)	F�TP��?'?�?K7��mment T�BD�?u7 >)�ETHERNE�T�?f�!OHOC�Ethernet� �figura��/D�1DCSVR�F�?�?�?�OQ1%��@ verif�y all�O�M�,��EDIFF��O�O�OO_R0%�HdiffQ_W�!>�@CHGD1F_-_?_�_ f_�_S+P�Y2�_�_�_Xo� �_ooGD�3No5oGo�o �no�fUPDA�TES."pi�FRS:\ a}�DUpdates� ListafP�SRBWLD.C	M�hLr�c��PS_ROBOW�EL�?<�aHADOW�o�o�of�Q3�Shadow Changesi�ޗ=�&�NO�TI�OA�S��O5NotificqB<���O�AJ?� nc��p���D��L� �󟂟���;�M�ܟ q� �����6�˯Z�� ~���%���I�دm�� ���2�ǿٿh����� !�3�¿W��{�
ψ� ��@���d���ߚ�/� ��S�e��ω�߭߿� N���r����=��� a��߅��&��J��� ������9�K���o� ���"�����X���|� #��G��k} �0��f�� �,U�y�� >�b�	/�-/� Q/c/��//�/:/�/ �/p/?�/)?;?�/_? �/�?�?$?�?H?�?�? ~?O�?7O�?DOmO�? �O O�O�OVO�OzO_�!_�OE_�Oi_{_�$�FILE_LpPR�[p��_P�����XMDONLY 1a�U~ZP 
 �
_ �_._oR_o;o__o �_�o�o$o�oHo�o�o ~o�o7I�om�o � ��V�z� !��E��i�{�
��� .�ÏՏd�������� *�S��w������<� џ`������+���O� a�🅯���8���߯~�ZVISBCK�X|�Q�S*.VD�|0���FR:\���ION\DATA�\�â��Vi�sion VD file\�j����� ̯ڿį�����4�ÿ X��|ώ�ϲ�A��� e�w�ߛ�0�B���f� �ϊ�ߛ���O���s� ���>���b���� ��'��������� ��'�L���p������ 5���Y���}���$�Z�MR2_GRP �1b�[�C4�  B� 	 ��Qk}h E�� �E�  F@ �F�5U�/
h L����M��J�k�K�v�H�,�Hk���?�  �/h 9�tQv8����6h�%�A��  3EBHeB)�a `�E@i/�g��h @UU�U�U��>�]��>П�;r�8	===E���<D�><��ɳ<�Ε�:��b�:/'79��W�9
@�8�8�9���T/�Q/�/eE7� E?p D�D��/�D�  D��  Cζ/9
_C�FG c�[T ��/?0?B?�N�O �Z
F�0x1 }0�RM_�CHKTYP  ��P� �P�P�P���1OM�0_MIN��0
���0�P]X�PSSB�#d�U�Pi�?	��3O$O�UTP_D�EF_OW�P
|�Y?AIRCOM�0�JO�$GENOV_RD_DO�6�RnxLTHR�6 d�E�d}D_ENBiO �}@RAVCGe��7� ��Fn�H E�� Ga� H�� H�?@Jh`�/O�?_�G_X_{ ���AOU�@kN� {NB{8���_y_�_�_�_/  C�� 	$o�X0YoilCOmB��AVbp~	�Y+O�@SMT�C�l�IZ �04d�$HoOSTC�"1m�o� 	
xM
{
:byeV���� �zu� ��$�GH���p	anonymousK�y������� ��	-�A�c �V�h�z������ ԟ����M�_�@�R� d�v���ˏݏ��� �7��*�<�N�`��� ��������̿�!�3� �&�8�J�\ϟ���ï կ׿��������"� 4�w�X�j�|ߎߠ��� ���������0�s� �ϗϩϫߜ������� �����K�,�>�P�b� ��s��ߪ��������� G�Y�k�L�p�� ������  $6YZ��~�� ��	�-? /S uB/h/z/�/�/��/ �/�/�/
?-/_qR? d?v?�?�?��// ?�?I/*O<ONO`OrO �/�O�O�O�O�OO3? E?&_8_J_\_n_�g�a�ENT 1n�i��  P!�O�_  �@�_�_�_o �_+o�_Ooo[o6o�o �olo�o�o�o�o�o 9�oo2�V� z�����5�� Y��}�@�v�����׏ ��������+��T� y�<���`�����埨� 	�̟ޟ?��c�&����J�QUICC0���p�!172.8.9.225�����1���ү3���2�4������!ROUTER��`�r�ӿ!PCJOGԿ���!192.�168.0.10�����CAMPRT,$� �!�1�K�2�RT��O�a��ψTNAME !�Z?!ROBO=����S_CFG 1m��Y ��Auto-sta�rted�4FTP�?[��?�O��O �߼������ߋO�(� :�L�o�]����������#��:4�F� X�9�l��P������� ��z�������#F� ��Yk}����?�=SM�65233)�
=_�,R dv�K�����  %��5/G/0Y/k/}/""q��? �?�?�/3?&?8? J?\?/�?�?�?�?�? �/m?�?O"O4OFOXO �/�/�/�/�?�O?�O �O__0_�?T_f_x_ �_�_�OA_�_�_�_o o,ooO�O�OEo�_�o �O�o�o�o�o�o( :L^�o��� ��� �CoUogoH� {�o�������Ə� ���� �2�U�׏U� z���������)� ;��O�q�R�d�v��� ��]���Я����)� ��<�N�`�r�������_ERR o�������PDUSIZW  3�^L��ȴ�>�WRD ?�"���  guest-��!�3�E�W�i�{���S�CDMNGRP �2p"�˰C��3��-�K��� 	P01.0�5 8�� ������> j  2��1�� � ����T���������������$���ϿQ�<�u��`�������  �  
���N(�P,�(�����Q����������l�� 8�#{�d�����|"ߙ�_GROU��Uq������	�����4S�QUPD � �ȵX��T�Y�����TT�P_AUTH 1�r�� <!i?Pendan�����8�g�!KAREL:*�����KC-�=�O�%��VISION SCETb�����!�� ����"� ��_�6H�l~��CTRL s������3���FFF9�E3��FRS�:DEFAULT�FANUC� Web Server����	�� �}��������WR_CONFI�G t�� ���IDL_CP�U_PC*3�B���I  BH/%M�IN:,��M%GNR_IO�����Ƿ1 �NPT_SIM_�DO&�+STA�L_SCRN& ���*TPMODN�TOL�'�+bRT�Y�(I!�&����EN�B�'��-$OLN/K 1u���Q?�c?u?�?�?�?�?52M�ASTE~ ��52SLAVE v��|34��O_CFG�?�IUO��OBCY�CLE>OD$_A�SG 1w����
 �?�O�O�O�O�O �O__1_C_U_g_y_��_�;tBNUM�zĹ
BIPCH[O���@RTRY_CN*�"ĺB�!��P1�ȵ B;@B�x�>�Jo�1 SD�T_ISOLC � ��f��$J2/3_DS4�:�~�`OBPROC?n�%JOG^�1y�;���d8�#?��[�o�_?؟֟O|QNs��V����-�~o�h�`�Y A�_�bPOSR�E�o�&KANJI�_�0���/k�+�MO�N zg��2�y �Ϗ����Ҿ)�0c{,�9�T���e�_LY �R�_k�EYLOGGIN@�����ȵ�$�LANGUAGE� k2$ ,㑱�LG1b|�2�K��3�x�������O � '0,��W �
q�3��MC:\RSC�H\00\��L�N_DISP �}�?f�MKm�O�C�"@"Dzh#�A��OGBOOK ~K��w���w�w���X���-�?�Q��c�u���11����	���h�޿�����ॐ_BUFF 1@=��� )�����E�a�sϠ� �ϩ���������� B�9�K�]�oߜߓߥ���ߜ��DCS }�� =��͗� ֿM�l:�L�^�p����IO 1�K No��������� ������%�9�I�[� m������������������!3EY��Ex TMlnd��� ���0BT fx��������//���SEVt`}��TYPln���/�/�/)-P�R�S�P���bFL 31���`��?�,?>?P?b?t?�?�/T�P��loq"��NG�NAM�d��Ւ��UPSu�GI�U\�e}�1_LOAD�`�G %}�%D?F_MOTN$�FO�ݠMAXUALR�M�Wk�X\@�1_P�R�T`ԣ��Z@Cx��ꩦ��OV�9ż�C�`P 2��Kk �9�	q!P]  ��OQ�R 9_$_6_o_�]_�_�_ �_�_�_�_�_oo@o Ro5ovoao�o}o�o�o �o�o�o*N9 rUg����� ��&��J�-�?��� k�����ȏڏ����� "���X�C�|�g��� ����֟����ݟ�0� �T�?�x���m����� ү��ǯ��,��P��b�E���q���SGD_LDXDISA�0��;��MEMO_A�P�0E ?�;
 j ����*��<�N�`�rτ�Z@IS�C 1��; � ����T�A���ϛ�$���Hߙ�C_MST�R �B-g�SC/D 1����<߶� 8���������"��� X�C�|�g������ �������	�B�-�f� Q���u����������� ��,<bM� q������� (L7p[� �����/�6/ !/Z/E/W/�/{/�/�/ �/�/�/�/?2??V?�A?z?e?�?�?�?X�MKCFG �v���O�CLTARM_*�2��G�B P�2��@>OFD{@METP�U�C�@��~�ND>�@ADCOL`E�@�kNCMNT�O tEo� �v��N5C�.A�O�DtEPOSC�F�G�NPRPMl�OYST@1���� 4@��<#�
oQ�1oU_�Wk_�_ �_�_�_�_�_o�_o Oo1oCo�ogoyo�o�o�o�o�atASING_CHK  �O�$MODAQC���?���>+uDEV �	��	MC:>_|HSIZEѽ����+uTASK �%��%$1234?56789 ��u�)wTRIG 1�
��l#E%��)����0S�6�%C�vYP�q>��At*sEM_IN�F 1�#G� `)AT?&FV0E0`�׍�)��E0V1&�A3&B1&D2�&S0&C1S0}=ƍ)ATZ׏+��H/�W��K���A����j�ӟ����	� ��.����� ��;����Я⯕�� ��*�<�#�`��%��� I�[�m�޿鯣��K� 8����n�)ϒ�y϶� ��{��ϟ���ÿտF� ��jߡ�{ߠ�S���� �����������T�� �+ߜ��a���	��� ���,���P�7�t��� 9��]�o����� (:q�^��=����XNITO�R�@G ?s{  � 	EXEC�1�32%3%4�%5%�p'7%8
%9�3 ��$ �0�<�H�T �`�l�x����2�2�2�2��2�2�2�2��2�2�3�3�30+qR_GRP_SV 1���� (�a��\���*X>�<����A���#c�>��~Z}�q_D�{�~�1PL_NA_ME !#E0��!Defau�lt Perso�nality (�from FD)� �4RR2�! 1��L68L@y�1P
d d�? v?�?�?�?�?�?�?�? OO*O<ONO`OrO�O@�O�O�O�O�OJx2e? _ _2_D_V_h_z_�_�_�_r<�O�_�_�_ o"o4oFoXojo|o�oH�o�i�V�_�n
�o�oNtP�o*<N` r������� ��&�8�n��� ������ȏڏ���� "�4�F�X�j�|�K�]� ��ğ֟�����0� B�T�f�x����������Ү FnH F�� G=��'�   �����"d���0�B�&�d�r� �׭Ҫ\�������ݿ� ͸��� � �0�6�T�vϿ ��|��ͰA�  �� ˿��Ǹ]0���ƿ3� ¿W�B�{ߍ�x߱�B5�K3�9^0`�!?0 � �0~�� @D�  ��?����?� ��!A�����$��(�;�	l�	 ���p��V� ]0M� � �/ � �l�r� �K(��K(��K ��J�n��J�^J&ǂ��2������� @�Y�,@Cz@I�@���������N����f����_�I����SѬ�Ä���  <��% �3�������!?s�8y�
�/�!��x����T� ܀��������}���    �������  ����������	�'� � 0�I� �  y�����:�ÈT?È=���l��	�(|�����ѦD���ψ��N@0�  '����@2��@���Y@!����@)��}C@0C��\CI��CM�CQ�� ���ģ�%%����� ����B���@0��l1@� ��!Dz����V�//+/Q/���� �H@q)q6�%  ��+���� p�!?�ff0���/�/V/ ���/;��8� !?/:��D4�� \6Pf8�)c�\�\��?Lv �$���;�Cd;�pf�<߈<��.<p��<�?L:D��ݧA���d��|��?fff?��?&@��@��� B�N�@T� ,E�	��	A���dO �O�7H��/�O�O�O �O _�O$__H_Z_E_~_�MEF�m_�_ i_�_UO�_yI�_2o�X�C��E��"Gd G;ML!o�omo �o�o�o�o�o�o�o$ H��iww9��_ �o�U��*�<�ڪ����/�6�������ď��菎�A�A�����C؏=�ԏ��X��񨑟,���>��  �P��"@�z<��E� C���s��x�؄�(������/�B�/B"��}A��#A���9@�dZ?v�ȴ,��~���<)�+� =��G��j���q����
AC
=�C��������� ��p�C�c�¥�B�=���ff��{,�I����HD-�H�d@�I�^�F8$ �D;ޓܪ�̠J�j��I�G?�FP<����QpJnPH��?�I�q�F.� D��Ɵg�R� ��v��������п	� ��-��Q�<�Nχ�r� �ϖ��Ϻ������)� �M�8�q�\ߕ߀߹� �߶��������7�"� [�F�k��|����� ������!���W�B� {�f������������� ��A,eP� t������ +;aL�p�����(����3�:��1��%�3��V��/"��(/:/�!4M��xT/f/F1�=Ӏ/��/4Ue'��T9�-�)�/�/?�/4?�"<]�P�2Pf>�q ��?��?�?�?�?�9���(�?�?/OO0?OeOPO�QB�hOzO �O�O�O�O�O�?t.__R_@[/X_b_�_`�_�_�_�_�Q{f�_��_o
o@o.odorj  2 FnH"��F��"�G=��B# ��C9)��@|��@��o �q�o{E��� F��`�H C�����oA`�m�kE�0wGa�O����{?ސ�q ��\d  zq: `�
 �!� 3�E�W�i�{��������ÏՏ�������q ���P+�~Y���$MSKCFMA�P  �%� ^f�q�qp��D�ONREL  �X5[��0D�E�XCFENB��
8Y����FNC�����JOGOVLIMҍ�d����dD�KE�Y�����_P�AN����D�RU�N���>�SFSPDTYw0�������SIGN����T1�MOT럜�D�_�CE_GRP 1-��%[�\�O� �O�&��d�Q��u� ,�j���b�Ͽ��Ŀ� ��)�;��_�σϕ� LϹ�pϲ��Ϧ��%� �I� �m��fߣ�Ov�D�QZ_EDIT���U��TCOM_�CFG 1�Q������"�
��_A�RC_��X5ؙT�_MN_MODE���縙UAP_�CPLF４NOCHECK ?Q� W5�H���� ������'�9�K�]��o�����������v�N�O_WAIT_L؉��׾�NT����Q��{_ERR�ȡ2�Q��1�  ��t���H*������`�OI�Px� ���������A�/����%p��w��Av���I8�?0|4��pd�BPARAMJ�.Q����߶��8so� =�`345678901� / *�?/Q/-/]/�/��/u/�/�/�+�7��?<�7?��UM_?RSPACEN�'2�$�p?z4�$ODR�DSPE㌦��OF�FSET_CAR8�Ќ�6DIS�?�2�PEN_FILE��0�$��֌1PTION_IO
�=�@�M_PRG %�\:%$*IO[N�3W�ORK �Χ�� ���F7��B�h�� ��d�@(7�A	 ��x�A5���c��0RG_D?SBL  \5����|_�1RIEN�TTO��9�C���pZ��a�0UT_S/IM_DGX�+���0V�0LCT ��%�ҟDx=gT_P�EXh��?�TRAT�h� d���T�0UOP �u^�Ӡ��oo�_:oHi�$��2ǣ�L68�L@�_S
d d'?�o�o�o�o�o �o�o1CUg y�������I2~o'�9�K�]�o�@��������ɏ9�<� ���)�;�M�_�q� ��������H�j3� H1`��XRP�C� U�g�y���������ӯ ���	��-�?�Q� � 2���������Ͽ�� ��)�;�M�_�qσ� ��d�v��������� %�7�I�[�m�ߑߣ��������X���'��*��S�H�Z�?� }������&?�������������+� I�O�m����?@����>� A�  ���� ������M8q \����z�d`�O�P1�k�o��sd`�R�0 ��D$@ @D�  DD:?QD	���U�  ;�	l�1	 ��p�s& ' j� � � � ���� H<z�H<W�H3k7�G�CG���G9|+c	�H
���� CC9P/9P4�9S;Q9/�#�9 � ��  1!�H>7 3����/1/�C/�BY�����XQ�^�H�<Pq/ ܩ/�"2�#��3�.�  _  �0�� o�  0�6��/?�%	'� �� M2I� ��  ���
=����q?�;�#&�(�3�/�'�A�?4;�B��?�'NEPO C 'VP3D�b CEP_C��\Cf Cj �Cn/@OROߑ  �����D%%���� ��'B���FEP�E˜#@XP�E5z�_�s/8_#_H_n_�"�� �H]2�Y�A6�U  �C�H�A��0p�Q?�ff0���_�_s_ ��o(k�18�0>oLj-�!ad�'�0yfP�h�Y�yy�3?L�0�T�!�;�Cd;�pf�<߈<��.<p��<�?ijD��WA�Eل1d�3|1��?fff?�@�?&+p�$@���=r�N�@T� IuՉ��&q-�0!� �we o��� ���A�,�e�w�b� ������я����l�А�O��CE����2Gd G; �|>�����ß���ҟ ����A�,�e��� ��V����د6���r� #�5�G�Y��Z� �_ �f�������̿�
�&A @A�@%���5��C��Z���/i�?Ƀ؈Ϗ��ϳ�UģP��2]!YNE�� CU%�̣�Ŀ8����E�@I�!t��B�/B"�}�A��#A��9@�dZ?vȖ+�~��~��<�)�+� =�G��(߇Ԁ�q����
AC
=C������녡� ���p�Cc��¥�B=����ff��{��I���HD�-�H�d@I��^�F8$ D;����ڭ̠Jj���I�G��πFP<��Qp�JnPH�?��I�q�F.� D��E�τ�o��� ���������&��J� 5�n�Y�k��������� ������ F1j U�y����� �0T?xc �������/ />/)/;/t/_/�/�/ �/�/�/�/�/??:? %?^?I?�?m?�?�?�? �?�? O�?$OOHO3O XO~OiO�O�O�O�O�Oz��(}���3:�O�a��)U�E3�Vq�_+_9R�E_<W_t�4M��q_�_�t��=ӝ_�_4Ue'��T9�] �Y	o�_-ooQo?lz�%P�bP�n�����o��O�o�o�o�i���(L7\�mt�B����� ����o��K�9�o�]�/u������ŏ�ُ�{f��9��'�]�K�����  2� FnH��F�-Щ�G=��B@P!�F.�C9F��p��@2����	��C�E�� �F����H C� ��S�b������ ����¯ԯ��?���*��y�C�C�|�uC�}�
 ۯ >�P�b�t��������� ο����(ϧ��� ��m[�~Y���$PARAM_MENU ?�U��  �DEFPU�LSE4�	WAITTMOUT���RCV�� �SHELL_WR�K.$CUR_S�TYL����OsPT���PTB�����C��R_DECSN��teG�A�S�e� �߉ߛ߭������������+�=�f�a�SS�REL_ID  ��U�a�u�USE�_PROG %�p�%b���v�CCR����ax���_HO�ST !p�!�����T�`��8�����:�t���_TI�ME����a�GDEBUG��p�v��GINP_FLM3SK����TR����WPGA�� ��{��CH����TYPEm�y�a�[� �����! JEWi���� ����"////A/ j/e/w/�/�/�/�/�/��/�/??B?��WO�RD ?	p�
 �	RS��s�PNSu��~2J9O�rTE[��?COLu>8�?>�L�� �P��p����TRACECToL 1��Uz�w �` �������1LFDT �Q��U^@#@D� � sc01A kE{O�O�O �O�O�O�O�O__/_ A_S_e_w_�_�_�_�_ �_�_�_oo+o=oOo aoso�o�o�o�o�o�o �o'9K]o �������� �#�5�G�Y�k�}��� ����ŏ׏����� 1�C�U�g�y������� ��ӟ���	��-�?� Q�c�u�����gI���� ӯ���	��-�?�Q� c�u���������Ͽ� ���)�;�M�_�q� �ϕϧϹ�������� �%�7�I�[�m�ߑ� �ߵ����������!� 3�E�W�i�{���� ����������/�A� S�e�w����������� ����+=Oa s�������� '9K]o� �������/ #/5/G/Y/k/}/�/�/ �/�/�/�/�/??1? C?U?g?y?�?�?�?�? �?�?�?	OO-O?OQO cOuO�O�O�O�O�O�O �O__)_;_M___q_ �_�_�_�_�_�_�_o o%o7oIo[omoo�o �o�o�o�o�o�o� EWi{��� ������/�A� S�e�w���������я �����+�=�O�a� s���������͟ߟ� ��'�9�K�]�o��� ������ɯۯ���� #�5�G�Y�k�}����� ��ſ׿�����1� C�U�g�yϋϝϯ��� ������	��-�?�Q��c��$PGTRA�CELEN  �b�  ���a��w�_UP �����љ�В���w�_�CFG ������a������������׉���DEFSPD ����`щ��w�IN~��TRL ������8�F�PE_C�ONFI�Ш��O������WLID�ө��	��LLB 1���� t�?B�  B4��� ��� ����� 88�?�0�K�0�G�i�k�}� ������������5Ak��� ��2��	�?~��GRP 1����lb�A�  ��333a�A���D�@ D�� �D@ A@�Ta�d+������� 	='����#´#��B 9!�///O/9/s/
?��?����/�/��.�/ =o=	7L�/?�/?P? ;?t?_?�/�?�??�?<�?�?  DzC Oa�
OHO�?XO~OiO �O�O�O�O�O�O_�O�_D_/_h_S_�_�Z!�a�
V7.10�beta1�� �Ax���R�y�y�Q?���Qo>�\)�QB0����PA��SBp���QA�9Sy�b
a�S �_2oDoVoho��Ap���"���o��o�o�o�Ҹө�KNOW_M  �|�֦�SV ���/���5O8 J\u_�k}��Ҕ���M]�z�Д��R	��%%��"��|���G� ��u��P@��a�]�a�q�m��`��MR]��}��&%O�P��$ӏ�KST]1� 1���
 4 ��vi�Q:��"�4�F� w�j�|�������ğ	� ���?��0�u�T�f� ���������ү���2� �a��<K��^35�G�Y�k���4���������5 ۿ�����6.�@�R�d��7�ϓϥϷς�8������
��M_AD  �����OVLD  ���G�PAR?NUM  ���߾��T_SCHy� ���
�����0�U�PD��������_CMP_�p|�pp�'�e��ER_C;HK�����j�⌝��RS��oW_#MO{���_��տ_RES_G�� � o����������� ����2%VI@zm`�R�4�\�l� �Q������S�ڰ �S�-�9X] S��x��S���� ��S�&��//S�V 1���a�q�@c?\�THR_INR��~��r�e�d�&MASS�/ �Z�'MN�/�#MO�N_QUEUE C���f"��a��N��U��N�&��0�END1;�79EX1EF?75\�BEE0'?>3OPTIO$7D��0PROGRAM7 %�*%0T/���2TASK_I�{ԍ>OCFG ��/���?"@DAT5A�s�+K��"�2��O�O�O�O�O�O �O_!_3_E_�Oi_{_x�_�_ROINFO�s�oM�
4[_�_
oo .o@oRodovo�o�o�o �o�o�o�o*<�N`�W�T�oL ؊	!A�K_%A�8+I�^�vENB|б}�)��v2��xG%A2���{ P(O8�4�F� C�e���z_EDIT �+O����DWER�FLg8|# �RGA�DJ ��:A����?"���!߆1��q�]��3?���A<@��v�%<�l�ӈ���q2Y�)��R	H0le��{"6�?
��A�F$�t$ܖ*z�/� **:�� "�����d�1�f�Ցd�[�_"U�#���3� E�s�i�{�������߯ կ�a���K�A�S� Ϳw���������9�� ��#��+ϥ�O�aϏ� �ϗ�߻�������� }�'�9�g�]�o��ߓ� ��������U����?� 5�G���k�}���� -����������C� U���y��������� ����q-[Qc ������I� 3);�_q���t&	>O@/Հ./ g/R$ݙ�/ߓU/�/Q/��/�/�PREF S�)�ՀՀ
߅?IORITY�72F}��MPDSP�1�яG7UTFǓކOoDUCT
A�:��/��OG��_T�G΀B���2TOE�NT 1� �(!AF_IN�Eq0OG!t�cpO6M!u�d%O^N!ic�mMOu��2XY"��v���X1)� ��O�OX0��O�O�E �O)__M_4_F_�_j_ �_�_�_�_�_o�_%o7o*�3"��=Y�yo��o��>��J�B�/�io�o��������AK�,  �0�q'9K]X5��7�pHANCE C�)��rrn{d�o��uyw	3�?"3ق��PORT_NUUMr3X0����_CARTREP�R0����SKSTAvq7 C�LGS @�ȍ��K�X0U�nothing �����̏܌������#��?k�TEMP �ɕ94����_�a_seiban �/���/��͟���ܟ � �9�$�]�H�Z��� ~�����ۯƯ���� 5� �Y�D�}�h����� ſ��¿����
�C� .�g�R�wϝψ��Ϭ� ����	���-��*�c� N߇�r߫ߖ��ߺ��� ���)��M�8�q�\����6�k�VERSI�P0�7�� d?isable�r<�SAVE ʕ:�	2600H8K44����,�!�0.�@�_Od� 	��{2$ /����X�e����	-;
��c�n� ��L��_�0 1˧K�� "����0URGEpB�0T6>5�WFF� DOr6�r�6W�0��"�WRUP_�DELAY ��;�R_HOT �%%&~1��+R_NORMALy�2���SEMI��"/�!QSKI%P���w�x��g/ ��/�/�/r-�5�/�' �/??(?�/L?:?\? �?�?�?l?�?�?�? O O�?"OHO6OlO~O�O VO�O�O�O�O�O_�O 2_ _V_h_z_@_�_�_��_�_�_�_���$R�BTIF?�RC_VTMOUT�B���`DCR�ϾE) �~!6�V�w C�r��A�.�/|'�j�!tb ��<��a�o�o�o �;�Cd;�pf�<߈<��.�>�]�>П���o��o'8}  8^p�������� ��$�1%RD�IO_TYPE � �.�EFP�OS1 1���  x����� Ώ���{����:�Տ 7�p����/���S�ܟ ���՟6�!�Z��� ~����=���دs��� �� ���D�V���=� ����¿]�濁�
ϥ� �@�ۿd�����#Ϭ� ��Y�kϥ����*��� N���r��oߨ�C��� g��ߋ��&������ n�Y��-��Q���u� �����4���X���|� ��)�;�u��������� ��B��?x� 7�[����� >)b��!�E ��{/�(/�L/ ^/�/E/�/�/�/e/ �/�/?�/?H?�/l? ?�?+?�?�?a?s?�? O�?2O�?VO�?zOO wO�OKO�OoO�O�O_ ._�O�O_v_a_�_5_ �_Y_�_}_�_o�_<o��_`o�_�o�o|�2 1ш�2oDo~o�o�o  &oD�ohe� 9�]��
��� ��d�O���#���G� Џk�͏���*�ŏN� �r���1�k�̟�� 🋟���8�ӟ5�n� 	���-���Q�گu��� ��ӯ4��X��|�� ��;���ֿq������ ��B�ݿ��;Ϝχ� ��[����ߣ��>� ��b��φ�!ߪ�E�W� iߣ����(���L��� p��m��A���e��� ���������l�W� ��+���O���s��� ��2��V��z' 9s����� @�=v�5� Y�}���</'/ `/��//�/C/�/�/ y/?�/&?�/J?�/�/ 	?C?�?�?�?c?�?�? O�?OFO�?jOO�O�)O�O�o�d3 1� �o_OqO�O)__M_SO q__�_0_�_�_f_�_ �_o�_7o�_�_�_0o �o|o�oPo�oto�o�o �o3�oW�o{� :L^����� A��e� �b���6��� Z��~������Ə � a�L��� ���D�͟h� ʟ���'�K��o� 
��.�h�ɯ���� ���5�Я2�k���� *���N�׿r�����п 1��U��y�ϝ�8� ����n��ϒ�߶�?� ������8ߙ߄߽�X� ��|����;���_� �߃���B�T�f�� ���%���I���m�� j���>���b����� ������iT�( �L�p��/ �S�w$6p ����/�=/� :/s//�/2/�/V/�/<�O�D4 1��O�/ �/�/V?A?z?�/�?9? �?]?�?�?�?O�?@O �?dO�?O#O]O�O�O �O}O_�O*_�O'_`_ �O�__�_C_�_g_y_ �_�_&ooJo�_no	o �o-o�o�oco�o�o �o4�o�o�o-�y �M�q���0� �T��x����7�I� [���������>�ُ b���_���3���W��� {������ß��^�I� �����A�ʯe�ǯ � ��$���H��l��� +�e�ƿ��꿅�ϩ� 2�Ϳ/�h�ό�'ϰ� K���oρϓ���.�� R���v�ߚ�5ߗ��� k��ߏ���<����� ��5����U���y� �����8���\���� ���?�Q�c������� "��F��jg� ;�_���/45 1�?�� �n���f�� �%/�I/�m//�/ ,/>/P/�/�/�/?�/ 3?�/W?�/T?�?(?�? L?�?p?�?�?�?�?�? SO>OwOO�O6O�OZO �O�O�O_�O=_�Oa_ �O_ _Z_�_�_�_z_ o�_'o�_$o]o�_�o o�o@o�odovo�o�o #G�ok�* ��`����1� ���*���v���J� ӏn������-�ȏQ� �u����4�F�X��� �ޟ���;�֟_��� \���0���T�ݯx�� ��������[�F��� ��>�ǿb�Ŀ����!� ��E��i���(�b� �Ϯ��ς�ߦ�/��� ,�e� ߉�$߭�H��� l�~ߐ���+��O��� s���2����h���������9�16 1�<����2����� ����������R ��v�5�Yk }�<�`� ���U�y/ �&/���/�/k/ �/?/�/c/�/�/�/"? �/F?�/j??�?)?;? M?�?�?�?O�?0O�? TO�?QO�O%O�OIO�O mO�O�O�O�O�OP_;_ t__�_3_�_W_�_�_ �_o�_:o�_^o�_o oWo�o�o�owo �o $�o!Z�o~� =�as�� �� D��h����'��� ]�揁�
���.�ɏۏ �'���s���G�Пk� �����*�şN��r� ���1�C�U����ۯ ���8�ӯ\���Y��� -���Q�ڿu������� ����X�C�|�Ϡ�;� ��_����ϕ�߹�B����f�L�^�7 1� i��%�_������� %���I���F���� >���b�������� E�0�i����(���L� ��������/��S �� L���l ���O�s �2�Vhz� / /9/�]/��// ~/�/R/�/v/�/�/#? �/�/�/?}?h?�?<? �?`?�?�?�?O�?CO �?gOO�O&O8OJO�O �O�O	_�O-_�OQ_�O N_�_"_�_F_�_j_�_ �_�_�_�_Mo8oqoo �o0o�oTo�o�o�o �o7�o[�oT ���t��!�� �W��{����:�Ï ^�p�������A�܏ e� ���$�����Z�� ~����+�Ɵ؟�$� ��p���D�ͯh�񯌯 �'�¯K��o�
���<yߋ�8 1ז�@� R���
���.�4�R�� v��sϬ�G���k��� ��߳������r�]� ��1ߺ�U���y���� ��8���\��߀��-� ?�y��������"��� F���C�|����;��� _�����������B- f�%�I�� �,�P�� I���i�� /�/L/�p//�/ //�/S/e/w/�/?�/ 6?�/Z?�/~??{?�? O?�?s?�?�? O�?�? �?OzOeO�O9O�O]O �O�O�O_�O@_�Od_ �O�_#_5_G_�_�_�_ o�_*o�_No�_Ko�o o�oCo�ogo�o�o�o �o�oJ5n	�- �Q�����4� �X����Q����� ֏q���������T� �x����7�������MASK 1�û������XN�O  ���M_OTE  3�����i�_CFG ��p�����PL_R�ANGl�g�t�PO�WER �õ�ݠ|�SM_DRY�PRG %p�%�m���TART ��ծ#�UME_�PRO�����_�EXEC_ENB�  d�x�GScPDX�������gTDB��ϺRM޿�ϸI_AIRPUR�� p�B�<�ٛ�MT_�TРn���OBOT_ISOLC1��8������9�z�NAME �p�n�ۙOB�_ORD_NUM� ?ը5��H844 �g��bҘ ����/(/��^/Ҧ/����PC_TIMoEOUT�� x�oS232��1�4��γ LTE�ACH PEND�ANPЅ��������l�j�Mai�ntenance_ Consg�����"��f�No Use���߮����0�B�T��h�NPO�2�RҤ�z��e�CH_L[���p���	���!OUD1:���R됏VAIL��R�����x�e�PACE1� 2�p�
 ��濫��{鋓�������9˺�8�?�%���%���4 IDu�������Y�� ����):!4� 8�Uu���� ��/�):/!/O/ q���U/���/  ?�/?6??K?m// �/�/�/c?�/�/�/�? O2O	OOi?{?�?�? �?_O�?�?�OGO_._ @_'_eOwO�O�O�O[_ �O�O�_o�_+_<o#o Qos_�_�_�_Wo�_�_ �o�o8Moo �o�o�o�o�o�o�D ��4��I�k}� ��a���돽���0�B��+�X�2a� s�������W�͏������4�U�<�j�o�3 ~�������Ɵt��� �<���Q�r�Y���o�4������ѯ㯑�� )�8�Y��nϏ�vϤ�o�5��ʿܿ� Ϯ� $�F�U�v�9ߋ߬ߓ���o�6�������� ��A�c�r��V��������o�7����(� :���^�����s���������o�8�!�3� E�W�{���������o�G ��/ m�
nu d  / ������/N l -S-L/�/p�d� z��/�/�/�/ ??&?/./@.1:n? �;�?�/�/(?�?�?O O*O<O2?D?V?h?�? �O�O�?�?HO__&_ 8_J_\_ROdOvO�O�O�_ ` @ p��U]/o�O�IAakU�_Rodoj_DjEowo �o�o�o�o�o%�o �o=ASe� ��	���3�E��@�+�]���a�o\
#o��o�_MODE � /
�S �"/㏙_�Z�o�H�����	��㟐�CWORK_AD��
�O4��R  �/< 1���_?INTVAL�a��%�R_OPTI[ONR� %����V_DATA_G�RP 2�uX:D�@PП��̟�˩ ͏���1��U�C�y� g�������ӿ����� �	�?�-�O�u�cϙ� �Ͻϫ���������� ;�)�_�M߃�qߧߕ� ���������%��I� 7�Y�[�m������ ��������E�3�i� W���{����������� ��/SAwe�����P�$S�AF_DO_PULS�Q�A��� CAN_TIM���E}�R ���Ƙ�Eqsy�֡��Yo�K�C կ�� ����l//%/�7/I/[/e��C"�2�$KKd�(�!"�!ѢIf)�P5�@�/�/�/���)�/ ��~4�_ �R  T0�!?^?p?�?~�9T D���? �?�?�?�? OO$O6O HOZOlO~O�O�O�O�O��OU�s��'p�O$_6_�I  �T;�o��WQo��p�M
�t���Di��[=Z0 � ��o�[Q[S C�_�_�_�_o o2o DoVohozo�o�o�o�o �o�o�o
.@R dv������ ���*�<�N�`�r��������?��я� ����+�=�O���r% {�������ß՟��� ��"�_���02�S wU�]n���������ȯ گ����"�4�F�X� j�|�������Ŀֿ� ����0�B�T�f�x� �ϜϮ���������� �,�>ߩ�b�t߆ߘ� �߼��������o�(� :�L�^�p����� #�Q�[����
��.� @�R�d�v��������� ������'9K ]o������ ��#5GYk�}������ �O�3�//1/C/U/ g/y/�/�/�/�/�/�/ �/	??-?;:�D?\q?{6��d�j?�@]	12345�678�Rh!B_!����B��V��?�?OO )O;OMO_OqOwA��O �O�O�O�O�O__*_ <_N_`_r_�_�_�_�_ �]�O�_ oo$o6oHo Zolo~o�o�o�o�o�o �o�o�_�_DVh z������� 
��.�@�R�d�#�� ������Џ���� *�<�N�`�r������� ��y�ޟ���&�8� J�\�n���������ȯ گ����ϟ4�F�X� j�|�������Ŀֿ� ����0�B�T�f�%� �ϜϮ���������� �,�>�P�b�t߆ߘ� �߼�{�������(� :�L�^�p�����@������ ����0 .�@�%���l�~����Cz  B\�_   ��2d4�� ��d1
~���  	�d2�2,�%7IX%p���Z��� ����%7 I[m���� ����!/3/E/W/ i/{/�/�/�/�/�/�/ �/??/?A?S?e?w?D�?�:Z�����<�4���`�$SCR_�GRP 1��� �� �� ��� ���	 �1��2
BD[��� �� I�7GDO2OkO������hBDE� DP�wC�GhK��ARC M�ate 120iC 67890��wM-�@A 8��M2IA�A��?
12345�D;F�2  ����>U�1{F�1HC�1�A"hAJ<ANY	?R�_�_�_�_�_�\�G�H��0�T�7�2  o/O0oVoho7F/��Co�o?o�o���l0Q,�o:DBǲ��r�2tAA��A  @���YuA@�Wpj ?�wrH��Dz�AF@ F�` �r��o����� B�-�f�Q���}Yq�r`������ďքB�� y�*��N�9�r�]�o� ����̟���۟�&�@��CTOF�k������h�����qYq>���̣�7G@Ypݯ����W\HC+�3����AnpC�V��o~e$c��W��� y���������ո��¿ P�(�%�7��I�v�b�SS��0EL�_DEFAULT�  m�����u�HOTS�TR�͐���MIP�OWERFL  �������WFD�O�� �� u�R�VENT 1����`�� L!�DUM_EIP�L�(��j!AF�_INE��Fߺ�!'FT�u�<ߙ�9!o�� ������!RPC_MAIN���غ��1���'VIS��ٻ �}�o!TPp�PUt��/�dl���!
PM�ON_PROXY��2�e�������+��f�a�!RDMO_SRVb�/�gP����!RT��0�h,����!
��M,�,��i��E!RLSgYNCFl	84>�!ROS߸��4��!
CE>��MTCOM�2��k�)!	�CO�NS*1�lu!}�WASRC|��2�md�!�U�SB�0�n�/!�STM��'/.�o �Y/��}/p�J/\/�/��/�/�/��ICE_�KL ?%� �(%SVCPR#G1�/::$52:???")03b?g?)04�?�?")05�?�?)06�?�?)07OO)0
TJOE<	9ROWK&4��O)1 ,?�O)1T?�O)1|?�O )1�?_)1�?G_)1�? o_)1O�_)1DO�_)1 lO�_Q1�OoQ1�O7o Q1�O_oQ1_�oQ15_ �oQ1]_�oQ1�_�oQ1 �_'Q1�_OQ1�_w y1%o�/	2)0?"0� ��1�/��S�>�w� b�������я������ ��=�(�a�L�s��� ������ߟʟ��'� 9�$�]�H���l����� ɯ��ۯ���#��G� 2�k�V�������ſ�� �Կ���1��C�g��Rϋ��*_DEV ���MC�:��t����GRP 2�՟�0�bx 	� 
 ,����ߟ� ��7��[�B�Tߑ�x� �ߜ����������3� E�,�i�P������� z���������A�S� :�w�^����������� ����+O��D �<����� �'9 ]D�� z�����/h 5/G/./k/R/�/v/�/ �/�/�/�/???C? *?g?y?`?�?�?�?�? */�?�?O-OOQO8O uO�OnO�O�O�O�O�O _�O)__M___F_�_ �?x_�_p_�_�_oo �_7oo[omoTo�oxo �o�o�o�o�o�o E�_i{b��� ������A�S� :�w�^�������я�� ���^+��O�a�H� ��l�������ߟƟ� ���9� �]�D����� z����������� 5�G�.�k�R������� ſ��������C�p*�<�yϟ�d ���	gϰϛ��Ͽ����ό�+�%�+�Pߌ����i��i�y߇� qߧߕ��߹�����=� "�e���O�=�s�a�� ��������3��'� �K�9�o�]������ ���������#G 5k�����[�W ���C�j �3������ �/]B/�/u/c/ �/�/�/�/�/�/5/? Y/�/M?;?q?_?�?�? �?�/�?�?�?�?�?O IO7OmO[O�O�?�O�? �O�O�O�O�O_E_3_ i_�O�_�OY_�_�_�_ �_�_�_oAo�_ho�_ 1o�o�o�o�o�o�o�o Iooo@osa� ����!�E� 9��I�o�]������� �ޏ������5�#� E�k�Y���я����� �ן���1��A�g� ����͟W������ӯ 	���-�o�T�f��?� ��������Ͽ�G� ,�k���_�M�o�qσ� �ϧ�����C���7� %�[�I�k�m�ߵ��� ��ߥ����3�!�W� E�g���ߴ��ߍ��� �����/��S���z� ��C���?������� ��+m�R���s �����E* i�]K�o�� ��/A�5/#/ Y/G/}/k/�/��/�/ �/�/�/�/1??U?C? y?�/�?�/i?�?�?�? �?�?-OOQO�?xO�? AO�O�O�O�O�O�O�O )_kOP_�O_�_q_�_ �_�_�_�_1_W_(og_ o[oIoomo�o�o�o 	o�o-o�o!�o1W E{i��o�� ����-�S�A�w� ����g�я����� ��)�O���v���?� ����͟���ߟ�W� <�N��'��o����� ɯ���/��S�ݯG� 5�W�Y�k�����ſ� �+�����C�1�S� U�gϝ�߿��ύ��� ���	�?�-�Oߥ��� ����u��߽������ �;�}�b��+��'� ����������U�:� y��m�[�������� ����-�Q���E3 iW�{��� )�A/eS ����y�u� //=/+/a/��/� Q/�/�/�/�/�/?? 9?{/`?�/)?�?�?�? �?�?�?�?OS?8Ow? OkOYO�O}O�O�O�O O?O_OO�OC_1_g_ U_�_y_�_�O�__�_ 	o�_o?o-ocoQo�o �_�o�_wo�o�o�o ;)_�o��oO �������7� y^��'�������� ُǏ��?�$�6��� �W���{�����՟� ��;�ş/��?�A�S� ��w����ԯ���� ��+��;�=�O���ǯ ���u�߿Ϳ��'� �7ύ�����ÿ]Ϸ� ����������#�e�J� ���}�ߍ߳ߡ��� ����=�"�a���U�C� y�g��������� 9���-��Q�?�u�c� ������������� )M;q���� a�]��% I�p�9��� ����!/cH/� /{/i/�/�/�/�/�/ �/;/ ?_/�/S?A?w? e?�?�?�??'?�?7? �?+OOOO=OsOaO�O �?�O�?�O�O�O_'_ _K_9_o_�O�_�O__ �_�_�_�_�_#ooGo �_no�_7o�o�o�o�o �o�o�oaoF�o yg�����' �����?�u�c� ��������#���� �'�)�;�q�_���׏ �������ݟ��#� %�7�m�����ӟ]�ǯ ���ٯ����u��� l���E�����ÿ��� տ�M�2�q���e��� uϛωϿϭ���%�
� I���=�+�a�O�qߗ� �߻�����!߫��� 9�'�]�K�m���ߺ� �߃��������5�#� Y������I�k�E��� ������1s�X�� !�y����� 	K0o�cQ� u����#/G �;/)/_/M/�/q/�/ �/�//�/??7? %?[?I??�/�?�/o? �?k?�?O�?3O!OWO �?~O�?GO�O�O�O�O �O_�O/_qOV_�O_ �_w_�_�_�_�_�_o I_.om_�_aoOo�oso �o�o�oo�o�o�o �o']K�o��o ������#� Y�G�}�����m�׏ ŏ������U��� |���E�����ӟ���� ��]���T���-��� u�����ϯ���5�� Y��M�߯]���q��� ��˿��1���%�� I�7�Y��mϣ���� 	ϓ�����!��E�3� U�{߽Ϣ���k����� ������A��h�z� 1�S�-�����������[�@����$S�ERV_MAILW  ����e��OUTPUTt����RV 2�v	�  �� (�xO���i�SAVE���g�TOP10 2}�� d �� ;M_q���� ���%7I [m����� ��/!/3/E/W/i/ {/�/�/�/�/�/�/�/`??/?	�YP���f�FZN_CFGw �	����.��o1GRP �2�y7�� ,B�   A�0.D;� B�0�  �B4.RB2�1��HELLr2!�	��������7"O>1K%RSR1O2O DO}OhO�O�O�O�O�O �O�O_
_C_._g_R_��_�_�^�  ��%�_�_�_�R�\�a. �_b`)ރ��R2. do�_��6HK 1��; o�o�o�o�o�o �o�o
3.@R{ v�������<?OMM ��?2���2FTOV_EN�Bt����HOW_?REG_UIR�g��IMIOFWDL���!��5A��*SYSTEM*. �V8.30340� ł11/9/2�020 A ����X�SNPX�_ASG_T �  0 $AD�DRESS  ���ZE�VAR�_NAM	�%$�MULTIPLY���PARAM��� � $TgIME���$��_ID�	$NU�M�D�T�CIMP�[�FRIFD�VE�RSION��G�T�ATU �$DI�SK�NFOD�MO�DBUS_ADR8[�����PORC�`��SSR�� �x ��NGLE���g�$DUMM�Y7�SGL�T�ASK   �&����T������S�TMTT0�PSE9GT2�BWD�h���E��SVCNT�_GP�� 8 �$PC�ER_�V�   	$�FB�Pm�SPCX��m�ΐVDX�R[��� �$D_ATA00�u����1��2��3��4���5��6��7��8���9��A��B��C"��D��2���F�� Ty���1Ω1۩1�U1��1�1�1�U1)�16�1C�1P�1]�1j�1w�ҀIȪ��2Ω2۩2�2���2�2�2�2�)�26�2C�2P�2�]�2j�2w�3��3���3Ω3۩3�3���3�3�3�3�)�36�3C�3P�3�]�3j�3w�4��4���4Ω4۩4�4���4�4�4�4�)�46�4C�4P�4�]�4j�4w�5��5���5Ω5۩5�5���5�5�5�5�)�56�5C�5P�5�]�5j�5w�6��6���6Ω6۩6�6���6�6�6�6�)�66�6C�6P�6�]�6j�6w�7��7���7Ω7۩7�7���7�7�7�7�)�76�7C�7P�7�]�7j�7w����S�PRM_UPD~ӑ  $4�q� 
����ӑ�ؐ$TORQU�E_CMD   �u�MOa_SP�EEjQ_CURsREo�nAXI� �mS�CART��_Ut��̒�YSLO� � ��������䏐��_�{�VALU�OP��$�#(=F�ID_L��K%�HIF*IN�$FILE_A�v$�c$M�t��SAR0�  h^� E_BLCK���"��>�(D_CPU�)���)��F#y/�$���_�=�R 	 � 7PWҐOT��)1;LA#�SR� .3�?184RUN_FL�GQ5-4U184WIT X5v1-4v185H2�D4x�084̑TBC2��
 � $O��X0IGu �0_FT�M1D��42D�TDUCX0AZ��2M����6�1�7TH��C��DxGR.0A��E�RVE�3?D�3?D3�O��0_AC@ �X -$jAL�EN�3wD�3j@EL�_RATI��$&�W_�F#1jAc$2�GMO�!>��C��ERTIA�o!�I�aj@�KDE�E��LoACEM�CC�CmV�@MA��F7UW7QTCV>\_QWTRQ^\UuZ���C0t��USt�J_��q��M�TF�J2'���E�QUvA2�P>�s��a�C@JKfVK��1'a�1'a`A`J0l<d+cJJ3cJJ;cAAL+ca`3ca`[fe4\e5C�PN1�\P�`Q[;P�L�@_��E��3CF� =`^GROU1 �����y�N�0CC��`R�EQUIR*B��E�BUZ�fA�V$T�@2#qg@v�1��4 \�ENA�BL	�$APP�RpCL�
$O�PEN`xCLOSEEozSE�y�E
�1..� �u M�0<P8PB�t_MGr!�p�C��� �x��9P�wB{RK�yNOLD�v>h�RTMO_�3�$��uJ"��PcdP 3cP;cPcP�cPa6P��S�b� �4>�5� r�B��1���1��PATH��ӁɃӁ�Hσ0�r(p�W�SCATr��ar�qINiBUCh�@��)�C��UM2�	Y�@+@�P9�O!EA�T��0T�`@T�PAYwLOA�J2L7OR_AN�1��L*0����������uR_F�2LSHR9DؑL�O��(�ٗF��F�ACRL_�!&��"�䇔4bH$ �$H��rG�FLEXcs:�1J�6 PMr�?��?>OPO� c�iE :vO�FP٧��O5aP�O�O�LF1�>�R��O�O�O�O_!_��E+_=_O_a_ s_�_�_�_�_Y�vĽW �Sdf����_�_ o�jT2'W�X�`�e Ŵ��e'� �*o<oNo ``deme[ee�o�o�ot�i�2J�d ��0`�o�o� 8ATk�q�PELٰ}1=�x�J(p#pJE �C3TR"�f�TNR9��wHAND_VB�c�0 �� $���F2�v	D#S�W�!�3�v� $$M���yv�q��@�q�����>��AR  ���vQ!5��}A�| 
�zA�{A�@��{� ��zD�{D�P�G@0��ST�w���y��N�DYW0^p�v!� H���k@ϗ�ϗꑎ� g������PX�a��j�s�|������� Ģ�� ��Ť�����qASYM$��^�p������_�0�.�A�+��-��K�]�o�����J���K�����˙x�_�VI��	(�s V_UNIC.$P�בJeG"uG"�K$� X$|&
��P�K�,�>�d�%�T�\��à2�0H+0Rr���!Lv�VrDI�sO48�2� �c `�O�I2AO�F�I1l�W�W3o�~0�0ܰ�  � � ��MEB��@r2�"YT0PT���ڀ�1�`�dAu���8�1�9T���a $DUM�MY1`A$PSm_i�RF+�  ڀ��6XpFLA�`Y�P��B�3$GLB_T��5*E�0Vqp�`��j�v1 XMp�w��ST±#pS�BR��M21_V�rT$SV_ERb��O� pC�CCLD@�pBAڰOL2� GLv EW� 4�`��1$YQ�ZQ�W�C`ԑ��As02�����AU�E ��N��@�$GIz�}$�A �@�C�@�� L�`V�}�$F�EVNEA�R��Np�F]Y��T�ANCp���JOG��A� ��$JOINT
Ѻ`�"޶@MSET� E WECU۱�S��'U��� �g�U��?�#pLOCK_FO���0oBGLVm�GLhTEST_XMcpN�QEMP�Pr+bBB�P$U���B2�#2#p�CQab��4�PQarACE�`S�r` $KAR�M>3TPDRA�@�d��QVEC��f�PI�UQaVaHE�PT�OOL2��cV1�R�E�`IS3���b6�s�f�ACH�P(pb�aO��3�429�2��`ISr  @$�RAIL_BOX�E
��@ROBO�"d?��AHOWW�ARO�Aq�0qROLM�2gu��
txr�Ѹ/pZ���O_F��!G �D�a� �^*�PR�`Oˢ!�R*�d�Q�p�0�COU�R	"XBMeYC���P_$PIP#fN����b/r�ax�Qa�p��CORDED�P��q�� ��OY0 # 7D )@OBu�G� �Pd�S��3(@S��I�wSYSS�ADRH�� �0TCH�S� M,0EN2�A�Q�_T������PV�WVAu1% �� �`�B5PRE�V_RT�$E�DIT�VSHW�R��\F$����A�	 D�0��;���$HEAD�� U����KE�A�0C�PSPDl�JMPzp�L5L�TR��F44&[�t���I,`5SH�C��NE�`Iង�TICK2�<M�}����HNRA'� @]�����t�_GqP�&v��STY��qLODA�㖒��m�_( t 
 �GƅS%$�T=\@S>�!$=!2��1EF0rFP�SQU�`x%�B!TERC�0�Q���S��)  Ph@�׹���g��a�`1O�0�3t�IZDQE�1PRE��1!�̯��pPU�1�_DYObR��XS�PK6�AXIP��sVaUR�ڳI�Hp�~����_�`��ET��P( bl�O�FP�A�4 ss�`���SR��*lѠ�������� ���#��1��A� R�c�R�s�RŃ�d�~� ��dŢ������ː́C��|����S}C,@ + h�@cDS��a�0SPC0&~�ATq��2������2ADDRESz�cB�SHIF�^H`_2CHH�z��IK@���TV�I�72,��h���� 
�+j
��V�qA���- \����O������<�C��򢵲����B<��TXSCR�EEU�.	0k�T�INA�CP��Tp�Q����� / T�� �@����Ag@��^���8^����RROL wP`��f���v��QUE��G0 �� ��@S�Aΐ�RSM�T�UN�EX��6F�� S_ �Cf�6V�i���6���C�RB��� 2/��UE�1=2�B���!�GMT� Li!�m�w@O�wBBL_rpW�0��2 �O�jO�ALE���GpTO�3RI;GH&BRD�D���CKGR�0NTE�X��OJWIDT�Hs1�u�"qA�a�%�I_�0H�� '3 8�!wP_T�����0R�@�Rsw�2�$� O�ѭ�4��$�GG U2 �R brq�LUM�u���ERV
��@� PaP�У�5{0�GEUR�&cF���Q)]�LP$M��E��C�)jSѠx�x�`w5u6
u7u8Z���3�P9P��6�a�QS���4�USR�D'6 <���0UR���RFOC�aPPR�Iαmp�!L TR�IP+qm�UN$0547	Pt�$05�Yq5%�Ia���� q8�  �G \�aT�p1��ѣ"OS�1��&R���#�a�9��O�C�N�"�$�IaUU�:�/�/�U�N�#OFF!`��;[��3On0 ٰtW5�4:�@GUNw��P�0B_SUB8�2p@��SRT� �a<��vQ�p �ORpN�5RAU��4T�9䶇�1_���= |����OWN� T�$SRC���r�Dx!`CE�MPFI*�*ё�ESP-����� �e*B�&�b�!B�n��> `10WO8�rT�COP:1$��� _^@�b�A,�q�EWA�C?a�A�@�C�A�C �VC�CH�? �qC?36MFB1���Q�VC4�Y`��@x# %rT���XdP^Ȕ�spC�pRUDRkIV���_V��uT̐fpD�MY_UBY�ZTV�����B���V�a�RP_�Sp�+��RL7�BMv$��DEY��cEX����EMU��1X7d[�US���p�o��G��PAC3INΑ}�RGMAad�wbF3wb3wb���ARaE����a�r7S�wb�pA R�@G�PP�r�`5VR� �pB !d�_���2	�BN��RECcSWo`_A$pa�8c�O!��QA��1s�E�UB��� �q5VHKG�C��Iz���.p��zsEA���w�@� 1u5U�MRCV��D ��FOS�M� Cs�	p�rX3�c�rREF�� �v�v�q p7��p  �z��z��{;��vpA_@@�zq��{��S�0/g�Sᡏ�髿d��E �$�=�ߠ) �UӠOU��b��ZS @�e2�2��$��R� �ΐB��2Ѻ�Kq�SUL6s�C�@CO:�� 3D)`�NT�CZ���BY��e�!e�$�L��S���S�����!��JTǤFt +��ǱT� ��CACH+�LO����*`�����@ܣC_LI[MI��FR%�Tj��'���$HO� 6B��COMMpSB�O�0 ]�Ԉ�I؄h@V�P�b��_SZ3dn���6����12����[`��&����AaM]P�FAI&�Gvt���AD��BMRyEׄ9�_SIZ��PH�`��FASY�NBUF�FVRTaDk�w�I�aOL��SD_@3��W3P�'ETUc�QNp[��ECCU�hVEM�`��۲&�VIRC���VTP�p{$��J�s�A�w�_DEL�A�cP�ƺ�KS��G��@9pCKLAS��3	ő_�F�ƀH$p"�S;��N��P/LEXEEI��B�/��4sFLK I  `]�^A��M���dwsP3S/�^@�bJ# ������#�#RS ORD@!� ��> 3 ނ�)�K��T\"����WwCb2V��g%L`�Qۑ6D4��\*b3UR4sp_R'�d� ��,a]��ծc�_od@&�{g��`B*�T�N'�SCO��*�C�  ad�"_f�"0�">�" K�"Y�J_\_nZ���� E\ AM�P�0� PSMf%M�p"%HADJT�/e��Bڒ� Np"q׬!�LIN]3q��XV�Rh$O\���T_O�VR� �ZAB�C�5P�bw�$��
�O�ZIPg%Qp"D/BGLV�CL�R ��纀ZMPCF��5R  r ���$\��QLNK�2
u�9M,a|�S �|q��^��CMCMi`C�C�C�ACtP_�  �$J:4D ��@QJ�V�4p$0�tO�UXW� ��UXE>a��E �[���	��u���T ����r��YK�D"0 Ut�"��^IGHbcFq�?( �K��>V � vG��$B$��@1e�B�҉�&GRV%�F� ���OVC�5�A7�w@(�`��
VBI���}D�TRACEB��V�1�SPHER>�P W , �3|I[�$SIM�Apz!� e#4P �e!0V&��qe!�m/!��%���/Kpb/t#�_UN�@_+fp&LCд�% �%�V M��ALIA�S ?e����%1�! ( he �!:?L?^?p?�?�66? �?�?�?�?�?	OO-O ?OQO�?uO�O�O�O�O hO�O�O__)_�OM_ __q_�_._�_�_�_�_ �_�_o%o7oIo[oo o�o�o�o�oro�o�o !3�oWi{� 8������� /�A�S�e�������� ��я|�����+�֏ <�a�s�����B���͟ ߟ����'�9�K�]� o��������ɯۯ�� ���#�5��Y�k�}� ����L�ſ׿���� ��1�C�U�g�y�$ϝ� ������~���	��-� ?���c�u߇ߙ߫�V� ����������;�M� _�q��.������� ����%�7�I���m� �������`������� !��EWi{& ������ /AS�w��� �j��//+/� O/a/s/�/0/�/�/�/ �/�/�/?'?9?K?]?�3�$SMON_�DEFPRO �����1� *SY�STEM*p:RECALL ?}�9� ( �}t�pdisc 0=�>172.8.9�.225:7864 4 *.*�;?13524 �2d?�O"O2L}tpc?onn 0 �?�?��?�O�O�O;G:co�py virt:�\output\�untitled�1.pc md:� over �09�1758336:?165386�O_�#_6L6�Bfrs:�orderfil�.dat�Dtmp_back\�? �O�_�_3_-�Bmdb:c@[_QMt_oo)o6<F1xFT:\�_cN@\B�_�o�o�o@B2FeaNo`o[Cyo
. �O�O�O�O���?C�
xyzrate 11 Qcu���*�=E�w�k4092 �������� =E�?Y�a�s���(� ;OML܏�2������ �vQ�c�u���*�=�O�968�����������P� a�s��� (�;�M�ݯ﯀����� ��ɟ[�m���"�5�<G�WB9756��� �ϗϩϼ�P� a�s� ��(�;�ML����2���ߣ�6H�l�88�022784:951580���#� 6_H_Z_R��ߎ��3� �_`�X�t���)�<o �o�o]���������o Q�c�`�y�
.A� S����������� ��u*=����� s��������^�� //&/���s�����/�/�/=�F�nE2�^@d/v/??+?>� ���'�/�/�?�?�?<߀NK\?n?�?O#O��7 FXN?�`�?�O�O��.�aO�8uO__*_r��3FOXHemp�\87`��O�_�_�_��+FV*.dZ_l\s_ oo(o;�M��S�_�_ �o�o�o��Rnaoso (�?M��o�o2����{�$SNPX�_ASG�������q� �P 0 '%�R[1]@1.Y1��y?���%� (��L�/�A���e��� ����܏��я���� H�+�l�O�a������� ؟����ߟ�2��<� h�K���o���¯��̯ ��ۯ����R�5�\� ��k��������ſ� ���<��1�r�U�|� �ϋ��ϯ������� 8��\�?�Qߒ�uߜ� �߫�������"��,� X�;�|�_�q���� ��������B�%�L� x�[������������ ��,!bEl �{������ (L/A�e� �����/�/ H/+/l/O/a/�/�/�/ �/�/�/�/�/2??<? h?K?�?o?�?�?�?�? �?�?O�?ORO5O\O �OkO�O�O�O�O�O�O _�O<__1_r_U_|_ �_�_�_�_�_o�_o 8oo\o?oQo�ouo�o��o�d�tPARAM� �u�q ��	��jP;t�Ap�h#t��pO�FT_KB_CF�G  s�u�sO�PIN_SIM  �{vu���p�pRVQSTP/_DSB^~r�|�x�`SR ay� � & S�OCKET�"���vTOP_ON_ERR  -�|Kx?�PTN �f�r�A;�RING_PRMI�� �`VCNT_�GP 2au&q�(px 	�̏p����ޏ��wVD��ROP 1�i'p� y�R�d�v������� ��П�����*�<� N�`�����������̯ ޯ���&�M�J�\� n���������ȿڿ� ��"�4�F�X�j�|� �Ϡϲ���������� �0�B�T�f�xߟߜ� ������������,� >�e�b�t����� �������+�(�:�L� ^�p������������� �� $6HZl ~�������  2DV}z� ������
// C/@/R/d/v/�/�/�/ �/�/�/	???*?<? N?`?r?�?�?�?�?�?��?�?OO&O0�PR?G_COUN�At��r�NuRBENBć�MEMwCAt�O_U�PD 1�{T  
;Or�O�O�O __(_:_c_^_p_�_ �_�_�_�_�_�_ oo ;o6oHoZo�o~o�o�o �o�o�o�o 2 [Vhz���� ���
�3�.�@�R� {�v�����Ï��Џ� ���*�S�N�`�r� ���������ޟ�� +�&�8�J�s�n����� ����ȯگ����"� K�F�X�j��������� ۿֿ���#��0�B��k�f�x�DL_INF�O 1�E9�@��	 �����������@�@��@�>�����.�
� ������A��/���%q��?w�Av���o���� Da���q~D�Q�?6���´�ߞ��O@YSDEBUG�\@�@��d�I��S�P_PASS\E�B?��LOG U���C����Θ�  ��A��UD1:\���_MPC�E��AH�� �Am�SAV �m�4�lL��S�SVd��TEM_TIME� 1	��@ �0����ă��_���$T1SVGUNYS�@]E'�E�r��ASK_OPTICON\@�E�A�A���_DI��xO��BC�2_GRP 2
�I=�����@�  �C�f�BCCF�G ���� l�]`]`ߕ ������� 7"[FX�|� �����/3// W/B/{/f/�/�/�/�/���,�/�/"?4?�/ ?j?U?�?y?�?���? ���0�? O�?$OOHO 6OlOZO|O~O�O�O�O �O�O_�O2_ _B_h_ V_�_z_�_�_�_�_�_ �_�_.oh� BoToro �o�oo�o�o�o�o�o &8\J�n �������"� �F�4�j�X�z����� ď���֏����� 0�f�T���@o����ҟ ���t���*�P�>� t�����f������ί ����(�^�L��� p�����ʿ��ڿ �� $��H�6�l�Z�|�~� ���ϴ��Ϡ���2� D�V���z�hߊ߰ߞ� ���������
�@�.� d�R�t�v������ �����*��:�`�N� ��r������������� ��&J �bt� ��4���� 4FX&|j�� �����//B/ 0/f/T/�/x/�/�/�/ �/�/?�/,??<?>? P?�?t?�?`�?�?�? OO�?:O(OJOpO^O �O�O�O�O�O�O _�O $__4_6_H_~_l_�_ �_�_�_�_�_�_ oo Do2ohoVo�ozo�o�o �o�o�o
�?"4R dv�o����� ����<�*�`�N� ��r�������ޏ̏� ��&��J�8�Z���n� ����ȟ���ڟ���� �F�4�j� ������ į֯T����
�0���T�>�r��$TBC�SG_GRP 2�>�� � �r� 
 ?�  ������ӿ ������-��Q�c��v�}���d0� ���?r�	 H�C�`�r���b�C�  B����Ȟ��>�ff�źƞH�������϶�\���H �h�BLcφ�B$дh�j߈ߎ߰�H�����ތ��@�@�� AƷ�f�y�D�V����������	��?33�3��2�	V3�.00��	m2;ia�	*T�L�pq�c�"����r����� ��l���_   ��B��X����u�J2}����5���CFG ->��� ��
��D��Go�o��
G��� ����5 Y DV�z���� ��/1//U/@/y/ d/�/�/�/�/�/�/�/ ????Q?����\?n? �?*?�?�?�?�?�?O �?1OOUOgOyO�OFO �O�O�O�O�O	_r�^� ._:�>_@_R_�_v_�_ �_�_�_�_�_o*oo No<oro`o�o�o�o�o �o�o�o8&\ Jl������ �����6�X�F�|� j�����ď��ԏ��� �܏.�0�B�x�f��� ����ҟ������� *�,�>�t�b������� ���ί���:�(� ^�L���p�������ܿ ʿ ��$��H�6�X� ~�(��ϨϺ�d����� �����D�2�h�Vߌ� �߰��߀�����
��� �@�R�d��t��� ������������ *�`�N���r������� ������&J8 n\~����� �"��:L
 �|������ �0/B/T//d/�/x/ �/�/�/�/�/?�/,? ?P?>?`?�?t?�?�? �?�?�?�?OOOLO :OpO^O�O�O�O�O�O �O�O_ _6_$_Z_H_ j_l_~_�_.�_�_�_ �_ oo0oVoDozoho �o�o�o�o�o�o�o 
@.Pv��T f������<� *�L�r�`��������� ޏ̏����8�&�\� J���n�������ڟȟ ���"��F�X�op� ��o>�į���֯� ���B�0�f�x���H� Z������ҿ��,� >���b�P�r�tφϼ� ���������(��8� ^�L߂�pߦߔ��߸� ������$��H�6�l� Z��~�������d� ���&�����D�V��� z�����������
 .��R@bdv� �����* N<^`r��� ���//$/J/8/ n/\/�/�/�/�/�/�/ �/?�/4?"?X?F?|? �?8��?�?�?t?�?�? OO.O0OBOxOfO�O �O�O�O�O�O�O__�>_(^  dPhS� hV|_hR�$T�BJOP_GRP� 20U�  ?�hVi	�R�S�\�8P���p���Q�U  � �� � ��RhS� @dP�R	 ��C� ff  �C�W�Q4b��|<f9o >�ff\a~<a=�ZC�`W���b�&`H&`!.g�o�gnѴW4e�\e`b�o ?a�d=߉7LC�noB��o#&`�`9u�o�c��33\uX2h�P<���C\vc@3?33@33|b}`��BL�wHqDa�l����u�Jh~�p<X��B$�d���?���C*p��C���Z`xy�x��k< �4�q`?]`C4.�Ϗ8R�d��daG�����{<g���]p@)&b`yap�c� z{4ep�V��������� �ʟ���(�� �N� �Z����������ޯ���d�hV0�4e	�V3.00�Som2ia�T*Z��TcQh�s� E��'E�i�F�V#F"wqF�>��FZ� F�v�RF�~MF����F���F���=F���F��ъF��3F����F�{G�
GdG�G#
���D��E'
�EMKE����E�ɑE�ۘ�E��E����F��F���F��F(���F5��FB���FO��F\���Fi��Fv���F��vF�u��<#�
<t���@Ť�r_X�j�M�hTn�@�U�S��SESTPARSA��\X�P�SHR��AB_LE 1�[��hS�ȃ� �0cɞǅ����gWoQ��	���
������hQ�������C���RDI�ϬQ��� �2�D�Vվ�O������ ����*���S�ߪS �������!�3�E� W�i�{����������� ����/A�]�� ���̂	k�}���M߀_�q߃ߕߧ���hN�UM  0U*�Q�PpP B�C�~��_CFG P��a@�PIMEBF_TT����S����VERAÔ�ޓR 1�[ �8e�hRcP! 3P�  � //$/ 6/H/Z/l/~/�/�/�/ �/�/�/�/? ?2?{? V?h?�?�?�?�?�?�? �>��?O�:0OBO TO.OxO�OdO�O�O�O �O�O�O_,__P_b_�8�_�_�_~_�_�_��_�_���_K�@����MI_CH�AN� � mcDOBGLV逡����p`ETHERA�D ?���`�n��?o�o�o��p`oROUT�!p
�!"t@|SNM�ASK�h��a255.~uF�|���F���OOLOFSg_DI��GT �i�ORQCTRL �p	��n��T �B�T�f�x������� ��ҏ�����,�>� P�b�r�����������PE_DETAI��h�zPGL_CONFIG Q�a��/cel�l/$CID$/grp1��3�E�W�i�{�1�	����ʯ ܯ� ���$�6�H�Z� l�~������ƿؿ� ������2�D�V�h�z� ��ϰ���������
� ��.�@�R�d�v߈�� )߾���������}��N�`�r��������턬��� )�;�M�_��߃����� ������l�%7 I[m������ ��z!3EW i������� ��///A/S/e/w/ /�/�/�/�/�/�/�/ ?+?=?O?a?s?�?? �?�?�?�?�?O�?'O 9OKO]OoO�OO�O�O��O�O�O�O_���User Vi�ew !�}}12�34567890 B_T_f_x_�_�_�T-`,��_��(Y25Y�O oo*o<oNo`o�_�_/R3�_�o�o�o�o�ogo)�^4�obt�������^5 Q�(�:�L�^�p�����^6�ʏ܏� � �$���E��^7��~� ������Ɵ؟7����^8m�2�D�V�h�z����럭��� lCamera3Z )����(�:�L�*�E�v�����@_��ƿ`ؿ�����  ̦ �Y�^�pςϔϦϸ� _����� �K�$�6�H�Z�l�~ߥ��̦�i� ������ ��$���H� Z�l�ߐ������� ��ߣ�Py��6�H�Z� l�~���7������#� �� 2DV��� *��������� ��"4F�j|� ���kͥ��Y/  /2/D/V/h/�/�/ �/��/�/�/
??.? ���l��/z?�?�?�? �?�?{/�?
OOg?@O ROdOvO�O�OA?�� � 1O�O�O
__._@_�? d_v_�_�O�_�_�_�_�_o�O�G9�_GoYo ko}o�o�oH_�o�o�o �_�o1CUgy
�	Υ0�o��� ����o2�D�V��o z�������ԏ{� Ӡիx�-�?�Q�c�u� ��.�����ϟ��� �)�;�M��ΥA�� ������ϯ�󯚟� )�;���_�q������� ��`��u��P���)� ;�M�_���ϕϧ�� ��������%�̿޵ ���q߃ߕߧ߹��� r�����^�7�I�[� m���8�޵�(��� ����%�7���[�m� �������������� ��޵���I[m ��J����6�!3EWi  	�������//(/:/L/^+   nv�/�/�/ �/�/�/ ??$?6?H? Z?l?~?�?�?�?�?�? �?�?O O2ODOVOhO zO�O�O�O�O�O�O�O 
__._@_R_d_v_�_��_�_�_�_b,  
� (  �( 	 �_oo:o (o^oLo�opo�o�o�o@�o�o �o$�Z~* ̸i{�  ������X 5�G�Y��}������� ŏ׏�����f�C� U�g�y��������ӟ �,�	��-�?�Q�c� ������������� ��)�;���_�q��� ʯ����˿ݿ��H� %�7�Iϐ�m�ϑϣ� ����� ����!�h� E�W�i�{ߍߟ����� ����.���/�A�S� e�߉��������� ����+�r��a�s� ������������� J�'9K��o�� �����X 5GYk}��� ���0//1/C/ U/g/��/�/�/��/ �/�/	??-?t/Q?c? u?�/�?�?�?�?�?�?:?p@ B"O4O�FOCG `��)�frh:\tpg�l\robots�\m20ia\a�rc_mate_}1�@c.xmlO �O�O�O�O�O__(_:_L_XX��X_}_�_ �_�_�_�_�_�_oo 1oCoZ_Toyo�o�o�o �o�o�o�o	-? VoPu����� ����)�;�RL� q���������ˏݏ� ��%�7�N�H�m�� ������ǟٟ���� !�3�J�D�i�{����� ��ïկ�����/� F�@�e�w��������� ѿ�����+�=�_H��1 Oj@8?8�?�=�|� =�xϚϜϮ������� �0��<�f�P�rߜ߀�ߨ��߼����&���$TPGL_OUTPUT "H1�H1 `� H�]�o������� �������#�5�G�Y� k�}����������������H�`���2345678901  2DVhz�>2 ������@9K]o�}� �������1/ C/U/g/y/�/#/�/�/ �/�/�/	?�/???Q? c?u?�??1?�?�?�? �?OO�?%OMO_OqO �O�O-O�O�O�O�O_ _�O�OI_[_m__�_ �_;_�_�_�_�_o!o �_/oWoio{o�o�o7o Io�o�o�o/�o =ew���E������+�� �} [�a�s���������̍�@b����h� ( 	 7�%�[� I��m���������ǟ ���!��E�3�i�W� y�����ï���կ� ����/�e�S����^�w���ѽ��� ��)�;���d�v� ϚϬϊ�����L��� ߺ�(�N�,�>߄ߖ�  ߺ���n������&� 8��D�n��^��� ������V��"���F� X�6�|�����z����� x�����0B��f x�����N `,�Pb@� ���p�/� /:/��p/�/$/�/ �/�/�/�/X/�/$?�/ 4?Z?8?J?�?�??�? �?z?�?O�?2ODO�? POzOOjO�O�O�O�O �ObO_._�OR_d_B_ �_�__�_�_�_�_o�o�_<oNoTb�$T�POFF_LIM� ���p��y��qibN_SVm`�  ӄjP_�MON #��)�d�p�p2Ӆia�STRTCHK �$��f^��bVTCOMPAT�h�q�fVWVAR �%�mAx�d ��o Y�p�b�ia_DEFPRO�G 3vb%S�OCKEp��m_DISPLAYt`��n�rINST_M�SK  �| ~�zINUSER��tLCK��{QU?ICKMENA��toSCRE`���~rtpsc�t��{���b��_��S�TziRACE_�CFG &�i�Atx`	bt
?�~܈HNL 2'�i}� �H{ nr4�F� X�j�|�������ĚޅITEM 2( �� �%$1234567890��  =<�7�I�Q�  !W�_�kp���bs�ů)�� ��_������^���y� ݯ����5�%�7�I�c� m�翑�=�c�u�ٿ�� ���!ϛ�E����)� ��5߱�����Yߧ�� ����A���e�w�@�� [�����ߧ��k� ��O��s��E�W��� c������}�'����� o�/������;S ����#�GY" }=�as��� �1�U/'/� �����_/	/�/ �/�/Q/?u/�/�/? �/i?�?�??�?)?;? M?�?O�?COUO�?aO �?�?�OO�O7O�O	_ mO_�O�Ol_�O�_�O �_�_�_3_�_W_i_{_ �_�_Koqo�o�_�oo o/o�o�oeo%7�o C�o�o��o����O�s�N�ڄS��)�S��  ϒS� �����y
 ��ݏď����UD1:\����e�R_GRP �1*��� 	 @�pY�k�U��� y�����ӟ��������͑�2��V�A�?�  q���m����� ǯ���ٯ�����E� 3�i�W���{���������	!����c�S�CB 2+o� \�Y�k�}Ϗϡϳ��������Y�V_CONFIG ,o��󁧏�M���OUT?PUT -o�>���Yߝ߯��� ������	��-�?�Q� c�u�;ъߝ������ ����	��-�?�Q�c� u�������������� );M_q�� ������ %7I[m�� �����/!/3/ E/W/i/{/��/�/�/ �/�/�/??/?A?S? e?w?�/�?�?�?�?�? �?OO+O=OOOaOsO �O�?�O�O�O�O�O_ _'_9_K_]_o_�_�O �_�_�_�_�_�_o#o 5oGoYoko}o�_�o�o �o�o�o�o1C Ugy�'�9Ո�� ����#�5�G�Y� k�}������oŏ׏� ����1�C�U�g�y� ��������ӟ���	� �-�?�Q�c�u����� ����ϯ����)� ;�M�_�q��������� ˿ݿ���%�7�I� [�m�ϑϣϴ����� �����!�3�E�W�i� {ߍߟ߱��������� ��/�A�S�e�w�� ������������ +�=�O�a�s������� ��������'9 K]o������ ���#5GY�k}����x�������/ �3/E/W/i/{/�/�/ �/�/�/�/�/?�/? A?S?e?w?�?�?�?�? �?�?�?OO*?=OOO aOsO�O�O�O�O�O�O �O__&O9_K_]_o_ �_�_�_�_�_�_�_�_ o"_5oGoYoko}o�o �o�o�o�o�o�o 0oCUgy��� ����	��,?� Q�c�u���������Ϗ ����(�;�M�_� q���������˟ݟ� ��%�6�I�[�m�� ������ǯٯ���� !�2�E�W�i�{����� ��ÿտ�����,���$TX_SCR�EEN 1.����}�ipnl/`�gen.htm,�ϑ��ϵ���$ Pa�nel setup��}�����0�B�T�f����ϝ߯� ��������n���?� Q�c�u����"��� ������)������� q�����������B��� f�%7I[m�� ��������t ��EWi{�� �:��////�A/�/�UALRM_MSG ?L��Y� Z//��/�/ �/�/�/�/??$?B?�H?y?l?�?�?�?u%S�EV  �-��6s"ECFG �0L�V�  �/�@�  A#A �  B�/�
  �?6�L�VOhOzO�O�O �O�O�O�O�O
_W�1�GRP 21	K; 0/�	 @Ob_�u I_BBL_N�OTE 2	JT��l6��Q�8�@uRDEF�PRO %�+ (%�?�_8��_o�_ 'ooKo6oooZo�o�o��o�o�o�ok\INU?SER  �]P_��oI_MENHI�ST 13	I  �('p ���(/SOFTPA�RT/GENLI�NK?curre�nt=menup�age,153,�17�����)�q�~381,23 �/�A�S��'��~71�����ӏ��qy+y��uedit�r?SOCKET��7� I�[���o������ǟ ٟ�z��!�3�E�W� i���������ïկ� v����/�A�S�e�w� �TEplq�����Ϳ߿ ���'�9�K�]�o� ��ϥϷ��������� �Ϡ�5�G�Y�k�}ߏ� ߳����������� 1�C�U�g�y���,� ��������	����?� Q�c�u����������� ����),�M_ q���6��� %7�[m ���D���/ !/3/�W/i/{/�/�/ �/�/R/�/�/??/? A?�/e?w?�?�?�?�? �����?OO+O=OOO R?sO�O�O�O�O�O\O �O__'_9_K_]_�O �_�_�_�_�_�_j_�_ o#o5oGoYo�_}o�o �o�o�o�o�oxo 1CUg�o��� ����?�?�-�?� Q�c�u�x������Ϗ �󏂏��)�;�M�_� q��������˟ݟ� ���%�7�I�[�m�� � ���ǯٯ���� ��3�E�W�i�{�������ÿտ��������$UI_PAN�EDATA 15����A��  	�}�/frh/cgt�p/widedev.stm�zό���ϰ���)prih��ϧ�}���"�4�F�X�j� )lߐ�w� �ߛ����������2� D�+�h�O�����������  w ������ ���#�5�G�Y���}� �ϡ�����������b� 1U<y�r �����	�-?&c�� D��C� ��������P !/��E/W/i/{/�/�/ /�/�/�/�/�/?/? ?S?:?w?^?�?�?�? �?�?�?Oz�=OOO aOsO�O�O�?�O./�O �O__'_9_K_�Oo_ V_�_z_�_�_�_�_�_ o#o
oGo.oko}odo �oO&O�o�o�o 1�oUg�O��� ���L	��-�?� &�c�J����������� ��ڏ���;��o�o ~��������˟ݟ0� �t%�7�I�[�m�� 柣�����ٯ����� ��3��W�>�{���t� ����տ�Z�l��/� A�S�e�w�ʿ����� ��������+ߒ�O� 6�s�Zߗߩߐ��ߴ� �����'��K�]�D� ����Ϸ��������� �d�5�G���k�}��� ������,����� C*gy`�� ��������}�,ew����)S�W��/"/ 4/F/X/j/��/u/�/ �/�/�/�/?�/0?B? )?f?M?�?�?�?�?Q������$UI_P�OSTYPE  ���� �	 �?#O�2QU�ICKMEN  �KO&O�0RE�STORE 16���  '��?X��O�C�OX�m�O�O__'_ 9_�O]_o_�_�_�_H_ �_�_�_�_o�Oo0o Bo�_}o�o�o�o�oho �o�o1C�og y���Zo��� R�-�?�Q�c���� ������Ϗr���� )�;����Z�l�ޏ�� ��˟ݟ����%�7� I�[�m��������ǯ ٯ�����
�|�E�W� i�{���0���ÿտ� ��Ϯ�/�A�S�e�w��1GSCREA@?�FMu1sc��@u2��3��4���5��6��7��8<���2USER����2��T����ks���U4�5�6�7��8��0NDO_CFG 7K<;��0PDATE ���������4B��_INFO� 18����RA0%}���Q�������� '�
�K�]�@��d�� ����������*L���OFFSET ;FM�Ë@ �b� t��������������� N�UL^�� �����&VO(�
L*�UFRA_ME  �d����RTOL_AB�RTp�ӈENB���GRP 1<��IRACz  A������	//�-/?&I/[/�@@U��iѠMSK  ���ӢNm%��%��/�_EV�N��$c�
6U�2�=I9hi��UEV�!td�:\event_�user\�/T0C�7Y?)�F�<L1S�PR1W7spot�weld�=!CA6�?�?�?�@�$!�/ h?&O[OGl�OJO8O �O�OnO�O�O�O_�O �O�Oe__�_4_F_|_ �_�_�_�_�_�_=o,o aooo�oBo�o�oxo��o�o'�o�j)6W�RK 2>@�88"�� y�� ��
��.�@��d� v�Q�������Џ⏽� ���<�N�)�_���~���$VCCMUҳ?\ݨ�MR�2�E8;<�"�	�j���~XC5G6 *����h֜ �5�i�A@�7 p? ȗ� ;[�e�Ȇ���ů�����^�9%A���ٯ*�� B���E��I�ѯ j�����]�����ֿ�� �����0χ��f�Q��cϜ�O����ϥ�ISIONTMOU?� ��ů�FU���U�(�� FR:\��\�u�A�?  ��� MC*�LOG�7�   UD1�*�EX[�E!' B@ ���Ҁo�r���o������d ��  =	 �1- n6  G-����Ҭ6,��<��1�=���:����n�P�TRAI�N����1�E!�Adt��͓G8; (�� :��S����������� -��1�?�Q�c�u���Й���T���_��REⲐH�����LEX�E��I8;�1-e���VMPHASE'  ���A����RTD_FILT�ER 2J8; ��R����� ��1C#�� t��������//��SHIFT6�"1K8=<���/p/3��O/u/�/�/ �/�/�/�/?�/?)? b?9?K?�?o?�?�?�?�	LIVE/S�NAP�3vsf�liv4�?�>�� SETU�0BmenuOO�?}O��OfB/%L����	|H{O�O��?�J� ��@-�AdB8
�����K�M�QR��S����	'-_�ME�0�ļ�/!M�OM �zWqW�AITDINEN�D����TOK C 噰\���_S�_�YTIM����
lG�_,m�_Ok�_/j��_/jo�XRELE�K_g���Q��֗Q_�ACT�0^h(q�X_N3� N��)r%�Ox_��rRDIS�0~�n�$XVR�B�O �$ZABCv͒1P�� ,��r��2g7ZIP�CQ����/�A�S��z�MPCF_G 1	R�J�0��w��a��MP�sS���<������8����v�4���?�  ������������m���Da���q~D�Q���?���\��*X�>�<���A����#c>��!~���"�4�;B�T� f�v�e�Ο����A�~2�6���´$� 6�>Ȇ�n�h�z�����ȫ�pt��T|��w�_YLINDqU|��  �e� ,(  *)�:���&�c�J���n� ���Ͽ �#��s�(��!�^� ���ϔϦ����e�K�  ���$��y�Z�l��{���2V�+q � ���������������٧�D��ז^�A����SPHERE 2W	�̾Ϛ�ߓ� �����<�O�*�<��� `������}������ ��I�[�8��\C�U�������pZZ�f ��f