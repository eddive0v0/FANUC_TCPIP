��   ��A��*SYST�EM*��V8.3�0340 11�/9/2020 A 	  ����CELL_G�RP_T   �� $'FRA�ME $M�OUNT_LOC�CCF_METH�OD  $C�PY_SRC_I�DX_PLATF?RM_OFSCt�DIM_ $BA{SE{ FSETC���AUX_OR�DER   ��XYZ_MAgP �� ��LENGTH�T�TCH_GP_M�~ a AUTORA�IL_  �$$�CLASS  O�����D���DVERSIO�N  ���/IRTU�AL-9LOO�R G��DD?8�?�������k,  1 <DwH8G���.��D@��82 ��-��Z�Z]/�o/�/S/�/�/�-_ ��/�/�/;�$MN�U>AP"�� 8 �'/�!I?�?m?? �?�?�?�?O�?O7O !OCOmOWOyO�O�O�O��O�O�O_�'5NU�M  ��	� �	�o%2TO{OL/?4 
E;zU�P���.Q13�P�Q��C�S_ )_+_�_�_o�_o=o 'oIoso]oo�o�o�o �o�o�o�o!K5@G�kdVIVy
WV6�