��   b�A��*SYST�EM*��V8.3�0340 11�/9/2020 A   ����CELLSE�T_T  � w$GI_ST�YSEL_P �7T  
7ISO:iRibDiTRA�R|��I_INI; �����bU9A�RTaRSRPNSS1Q23U4567y8Q
TROBQ?ACKSNO� �)�7�E� S�a�o�z�2 3 4 5* 6 7 8aw.n&GINm'D�&� �)%��)4%��)P%���)l%SN�{(O�U��!7� OPT�NA�73�73.:BP<;}a6.:C<;CK;�CaI_DECS�NA�3R�3�TR�Y1��4��4�PTHCN�8D�D>�INCYC@HG��KD�TASKOK�{D�{D�7:�E �U:�Ch6�E�J�6�C�6U�J�6O�;0U��:IATL0RHaRbH<aRBGSOLA�6�VbG�S�MAx��Vp��Tb@SEGq��T��T�@REQ �d�drG�:Mf�G�JO_HFAUL��Xd�dvgALE@� �g�c�g�cvgE� x�H�dvgNDBR�H<�dgRGAB�Xt�b�% LMLI�y@   �$TYPESIN�DEXS�$$C�LASS  ����lq�����apVERSION�ix  ���}qIRTUAALi{q'61�r���p��q�t+ U�P0 �xS�tyle Select 	  ����r�uReq. /�Echo���A�ck��Initiat�p�r�E
�^�m����ʠ�	��
��  ���������������χ�q)��O�ption biGt A<��p�B���C4�Decis��codY��Tr?yout mj�6��Path seg�h�ntin.8�I�g�ycX�:�Tas�k OK��?�Ma�nual optK.r�A���B����C� decs�n ��$�Robo�t interl�o7�@�\� iso)lQ�4�C��iM�@���ment<�)��������Ě}�stat�us=�	MH F�ault:����Aler�1�C��p@r7 1�z j�;��y���I�; LE_COMNT ?�y�   Չ�ѿ �����*�<�N�`� rυϖϨϺ������� ��&�9�J�\�n߀� �ߤ߶����������"�����U��Ђ��Ŵ�   ��ENAB  ��:��������������ꮵME�NU\��y��NAM�E ?%��(%$*R�זb��P���t� ��������������+ O:s^p�� ���� $ 6HZ�~��� ����/ /Y/D/ }/h/�/�/�/�/�/�/ �/?
?C?.?@?R?d? v?�?�?�?�?�?�?�? OM