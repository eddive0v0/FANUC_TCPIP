��   ��A��*SYST�EM*��V8.3�0340 11�/9/2020 Q   ���	�BIN_CF�G_T   X� 	$ENTRI�ES  $QW0FP?NG1FU1O2F2OPz �?CNETG  ��DNSS* �8 7 ABLE�D? $IFAC�E_NUM? $�DBG_LEVE�L�OM_NAM�E !� FT�P_CTRL.{ @� LOG_8	��CMO>$D�NLD_FILT�ER�SUBDI�RCAPdat��HO��NT.� 4� H�9AD�DRTYP� A H� NGTHOG�� �z +LS/� D $ROB�OTIG BPEEyR�� MASK@�MRU~OMGD�EVK� RCM�+ ;$��� ��QSIZ�NTIM$S?TATUS_�?�MAILSERV��  $PLANT�� <$LIN�<�$CLU��f<${TOcP$CC5&sFR5&JEC!}�ENB � �ALAR�B�TQP�w#�V8 S��_$VAR)M��ONt&��t&APPLt&PA� u%�s''POR �_T!["�ALERT5&2U�RL }�#A�TTAC[0ER�R_THRO�#UaS29�38� CH- ��[4MAX?WS�_1�y1MOiD�z1I� $y2� � (y1PWD � ; LAu00�N�Dq1TRY�6DE�LA�3z0��1ER�SIS�!�2�RO.�9CLK�8M� �Ο0XML+ �#SGwFRM�#TCP��OU�#PING_RE�5OP�!UF�#�[A�C�"u%_B_A�UZ�@��B�"CO�U!�UMMY1z�G2?�RDM*}� $DIS�I� J@Io/ 3 �$ARP�)_7IPFOW_�޳F_INFApD� �HO_� �INFO��TELs P~����� WOR�1�$ACCE� LV���RF�!�IC�E�0�Q �$AS ? ����Q��
��
�PV�1m@�W�  �5��QI0AL�_�QX'0 �X
���F��a���PBb;e��� #m��!�Qzo����$ETH_FL�TR  �Y.` U���������k��� #m2�kRSH�AR� 1#i G Pvo,8d XG|?�c�� �����B��f� )���M���q���䏧� �ˏ,��P��%��� I���m�Ο��򟵟� (��L��p�3���W� ��{�ɯ��կ6� ��Z��~�A�S���w� ؿ������ ����V� �z�=Ϟ�a��υϻπ�������@ߒgz _�L�11�mx!�1.{�0I��z�1|���255.��L�����@ey�2�߀���Ц߸�������3 �ߒ�o��0�B�T���4p������������5���_�� �2�D���6`���������Ȫ�������6A�MY�(MY���p��P�� Q� 8�< r������%7 �Pgy� J�����	//-/���Cew/b,�Q/��/�/�/�/�}�iRConnect: irc4�//alerts �/9?K?]?o?5�/�?@�?�?�?�?�?�0cP9a���?0OBO TOfOxO�O�O�O�O�O�O�O_�$�?3_�`("_[_�/_�_�_�_R����`a�i@�R>j�U�Q�Qt)�e�I DMZcan�$_TCPIP[b�m�i(`=aEL`���e�Q��`H!T�B�o�rj3/_tpdb/ m�vQ?!KCL�o�k�v_.��V!CRT��o�oF`�d!OCONSG�j�aOsmonL�d