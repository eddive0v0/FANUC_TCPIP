��  �A��*SYST�EM*��V8.3�0340 11�/9/2020 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA{RA�  ����ALRM_REwCOV�  � wALM"ENB���&ON&! MD�G/ 0 $?DEBUG1AI"�dR$3AO� TY�PE �9!_IF�� ` $E�NABL@$L�� P d�#U�%Kvx!MA�$LI"�
� OG�f �%�CAUSOd!PPINFOEQ/� �L A ��!�%/ H ��'�)EQUIP� 20NAM�r �72_OVR��$VERSI�3 ��!COUPL�ED� $!P{P_� CES0s!�o81s!Z3> �!� � $SO{FT�T_ID{2�TOTAL_EQfs $�0�0NO�2�U SPI_IND�E]�5X{2SCR�EEN_84o2SIGU0o?�;�0�PK_FI� �	$THKY-GP�ANE�4 � D_UMMY1dTD�d!_E4\A��A�R�!R�	 � �$TIT�!$I��N �Dd�Dd ��Ds@�D5�F6�F7*�F8�F9�G0�G�G@ZA�E�GrA�E�G1�G1�G1�G1�G �@~!SBN_CF>"�
 8F CNV_�J� ; �"�!_CM�NT�$FLA�GS]�CHEC��8 � ELLSE�TUP � 7$HOC0IO@� �%�SMACRO��RREPR�X� D�+�0��R{�UHM��PMN�B�! UTOBACKU��0 �)DoEVIC�CTI:0��� �0�#�/`B��S$INTERV�ALO#ISP_UsNI�o`_DO^f<7�iFR_F�0AINA���1+c��C_WA�d'a�jO�FF__0N�DEL�hL� _aAqQb�?Yap.C?��Y`A-E��#%sAT9B�d��AW{pT= $DB� g"z� S�$MO�0�B !kq� \v� VE~a$FN!��pd�_�t�rdT_MP1_F�u2�w�1_~c�r~b MyO� �cE D �[mp�a���RE�V�BIL0�!X�I� �R  �� OD�PT�/$NOnPM��I�b�/"_�� �m���H��0DpS� p E RD_�EL�cq$FSS�Bn&$CHKBD�_S�r�aAG G��"$SLOT_���2��� Vt�%𿃭3 +a_EDI�m   � ��"��PS�`84%�$EP�1�1$O�P�0�2qc�_OqKʂ� e0P_C� �c�+dR�U �PLACI4!�Q���( �ar�pM� <0$D������0pB�UOgB,�I�GALLOW�� (K�"82�0V�AR��@�2�sBLv�0OU7� ,yqȗ`7��PS�`�0M_�O]d���CFn�� X0GR`0���M]qNFLIx����0UIRE���$�wITCH�sA�X_N�PSs"CF�_LIM�t=�SPEED�!���P(��p�PJdV���u��u3z`�P6��ELBOF� �W��W��p� ���3P�� F B���1��r1堺�G� �� WARNM�`d܁�P����NST� CO�R-PbFLTR^۵TRAT�PT `>� $ACCQa�(N �r�pI�o"6��RT�P_S�r WCHG@I�Z�QT���1�IE�T��Y1݀�� x �i#�Qʂ�HDR�BJ; #C��2��3���4��5��6��7J��8��9V3l�M$��	3 @F TR�Q��$�V����C�FN�_U�pY�k�OpT <F �������#�I2q�LLEC7�>"MULTI�b�"��A!cj DET_��R  4F S�TY�"b�=*�)�2��o���pT �|� �&$L�>�+�0�P��u�!TO���E`�EXT�יၑ8B���"2����
�t k0F�RLƯ�r�q���� !D" �M��Qm� �蠋c�����"��G�1�ց�qM���P��! �����# L0	����P �pA��$JO�B,�ǰR�x@~�IG��$ d��������@ �K� l��弧o�s_M�0b% t���F� CNG0A�qBA� ��x��
�!v@��� ��z�0�P{`X�R·&ΰf��Pt�a�!��"J!�_)R��rCJ$�*(J)�D�%CHӽ��z@h�P�Z�@ '.�RO`�&�ס�IT�c�NOM_�`���S��pTE(�@�݉��P�ǭ��RA�0�2&"<�>�
$TFV w�MD3�T���`U(C1[�g�'�Hgb�s1q*E���\Ѕs�q�ŦgAŦsA�YNTt�q�P|pDEF�!)��G�PU8/@������AX��Ģ�ewTAI~cBUFņ����!sQ* � l�'�PI�)�P\7M[8Mh9� k6}F\7SIMQS)@�KEE�3PAT�Ѡ"�%"�"$#�"�L�64FIXsQ+ �ԭ�AdC_v�����23�CCIh��5PsCH�P�2ADD�6�,AE,AG,A!H�_�0�0_,@�foA)� ԀzFK� '�=$#�"�:�4E��, l���7@zpF�CE�C!F+H�S�EDIS�G�3�-z�P��MARG����r%�FAC
��rSLEW<�q�x;�,M��MCY.����pJB����
aC�W�v��U4��X/ ����CHNS_EMP��$GE g݀!_} ����pP�|!TC9f��y#a���Nd�W#%I��r<��<�J�R�И�SEGFRfoPIOj�ST`�gLIN׃�cPV����!�$0�����b�'��b�B��1` +`��	��a	`�� �a�Pܠ��At��Py�Q�SIZ���ltKvT`VsE pz�y�aRS%� ��uc@Q{k�|�`�xZ``Ld�| `�vCRCɥ��!����t�`%�p9a˭9b��MINQ��9a7��q�D�YCk�Cz��le����Lp ��EV���Fˁ_leF��N����Q(۶�X%+4,��#{0|!VSCA�} AY�=1)a/��2 �>�
/Ψ`_rU@� +�w][��i %�7��}R��3� �ߠ�߱���5ġR�HwANC��$LG��l�*1$�0ND�סAR�0NK�a�q��acm�ME�1��n��A0h�RA��m�AZ�����X%O`�FCAT���7`��S�P.
ADI�O��� ���pWP ������ⁱG��BMP�d�p�D&ah�AES�f@̓�W_P�BA�S���I9�4 � �I�T�C�SX@�w�5��	-$�1�T��?s�Cb�Ny`�aBP_H�EIGH71��WI�D�0�aVT�AC����!AQP0� �\��EXP+�L�@��C}U�0MMENU���6��TIT�1�	�%��aǱA1ERsRL���7 \��̉q��OR�D��_I�DG��QUN_O|d�L $SYS����4�ő�Iϡ	�E�VG#Ҍ�PXWO�����8.�$SK��*2�DBT(�T�RL��9 �� AqC`�u䈠IND� �DJ�4 _Z�*1XK�*�W�PL�A�R#WA.�tТSD�A���!�r@Y�UMM3Y9�ª�10����d���:	�A1PR�qw 
��POSr���; ��[$�$�q�PL��<��ߪS@��=�'�Cr�>4�'�ENE�@�T{�?S�S��R�ECOR.�@H� �O�@;$L��<$��62����0�`_q�b��_D9�W0ROx@�aT[���b��.�F��������P�Ac���bETURYN�V�MR��U� v��CR��EWM�b�mAGNAL� 72$�LA�e��=$=P�>$P٠= #?y�A<�C���@�DO�`����:�>��GO_AW ��MO�a)�o���C�SS_CNSTCY�@A L� ^�C`L' ID[^�2
2N��O����ـI�� B P�NPRB^rzCPI�POvI_BYȀR}�T�r��HN{DG.�C H��DQkSP�s*�SBLIO�F��0��LS�D��0N0�	3FB��FE���C��жE�DO&a-sO�MC`{P�4�C�rH��WFPrB=����SLA�P�F�bIN� �N3����G� $$���P]��v�� v�ޕ���!o�"�#ID�&L�&W��";$NTV*3"V9E 4��SKI��aHs�3�'2�b&aJ�x&aM�mdSAFE,d��'_SV��EXC�LU7ѻ���ON	L`�#YcL���4�ΤI_V8���PP+LYy�R��H[0'�3_M@�NPVR'FY_S�2MS�!O@��k6�1�~32�#Ot !5LS�E��#35�£1�`%�P��$��t5�%�g Hy��TA2МDP�� ҄S�G� I � 
$CURB�_�
� B�������#H��3F��UNM��DZD@���l�{IxA�X�J�F�EF��IM�J @F]Bk��pOTb�k�ԋѭ5��h�P�и@M� NI��!K��
RwPA!(T�DAY��LOAD�j��R�ӵ2 �E�F/�XILy�Ĉq}�OhPe�D�_RwTRQ�QM DF����P�r�S`�ThU 2L�`���Qkp�P���Q�QN 0�A��QA�t�R���DUtb���"�CAB�a�O�B�NS�QW`ID�`PW���U/q� �VjV_�P�P����DIAG�1�aP�� 1$Vb�HuT�l��u�t� �j���rR�p�DQ�tVE��Y@SW�ad�p7`q�d�U�PM�p�QOH�Uf�QPP�`�sIR���rB��Fb�S��q��q �@3r��-x ��-uj�#e�POwP�P���uR7QDWuMS���u�A�u�b�tLIFAEZ��C�p���rN�q �r�uxA�s�rI�xB�Cp���NC�Y���r�FLAW�y@O�V���vHE'ArSOUPPO2���rbS�_E�)E�_Xf�(h���s�Zp�Wp�p�`s���xA���XZ������qY2ˈC
�T������eN됕exAJJ� v_��q;���/���Q `[ CA�CHE��3�SIZ��v*��"j�N� UFFIo� �p��H�Ե3��6���M��R 8�@KEYoIMAG*�TM�င���D��q��O�CVIE�`�S �wP��Ll$@)#?G� 	��%���T�Pm�ST� !� �`!��@!�VP!��0!�EMAILy�1Q|��� _FAUL���U� �9��COU�z ��T��|aV<' $��zS�PC`;IT�#BUFF�)!PF�Oy�o�D�B���nC($����Ú�SAV�Ţ�`���`���|FP
�z���d�� _���"P_�OT�����P[0�Ѓ� B��AX��-�I���Wc�7�_G�s��YN_$q'�W�RDuY��U#rMb�T���F+�fP^@D�&�X�������g�C_��&�K��8�4B3���R��2�q��DSPl���PCy�IM� pÖ��#�Æ`UM�:���K0d�IPm#�q	�o�TH��=c�mPyT��p�HSDImƏABSCz$��o�V�� �Я�&�`ӀQNV�!GO�&ԑ�mƸ�	F�aаdR����,��SCxbk(�MER|4�FBCMP3��ET�1�Y��FUX�DU���\���%2CDf���z�u��R_NOAUT�  Z�P4 �"U��IUPS�C���C�1ϱב㍰���[H *�L  t�3���֚@�0�# �����A��VQ��1��扑��7��8��9P���p���1��1��U1��1��1��1��U1��1 �2�2�몥�2��2��2��2���2��2��2 �3J�3��3���3�ꨴ2����3��3��3� �4�}��EsXT�aQ\ < ���I簉���3�FDRxd]T��V�0���r�.�rREM�`F��r�OVMI�>AGT7ROVGDT�gMXvING�fNuaIND��r
�<�а$DG��:s�p��u�aD�VpR�IV���rGEA-RI�IO�eK7�tN�%(hQ�x0h `�>�sZ_MCMÀ�q�;�UR��^ ,<�1? �� s?� �a?�!�E�0�!ב����_�P}pP���`RI��դ$�aUP2_ g` VPģTD��@�3�#?@�!�'�%7�%wBACܲa T�hŢڠ�A);@OG.5�%�CT����IFI�q���x�:pC5PT|V����FMR2
�b �3LI��3#/5/�G/^|��u7_�D��R_�A�԰`M�|/-DGCLFuoDGDY_HLD�!��5�v��tz3�c��P�9 T�F9S]��d P� �B��0�а$EX_�A�H�A1kPl���@53[5V�G:�
ge ����SW�}O�vDEBUG4LWR�eGR� �U�ӷBKU��O1a� pPO�P�YoPع�BUoPMS�0OO,���QSM�0E�1��� _E f ��` �TE�RM�Ug�U}��O�RIe0�Qh�UFF �SM_80Ţ�P�i�Ug
�TA�ij'iUP�k� -��f$|�Ua`g$SEGfj�x@ELTOV�$wUSE��NFI"���bn �q+�d]dh$UFR02���a����	@OT�gU�TqA ��cNST`�PAT��?��bPTHJ ���E�:����bART+��e|�+��V��aREL<z9�S�HFT�a q.x_�SHI�M^���f �$`�xj)A�0OV9R��ǲSHI_p&D�U4� %�AYLO��AֱI�ѻ# qk�%�k�ERV���q� yz��g`<r4_0&�̥�_0RC�!9�AScYM	�9��aWJ�g��E�#*qV���aUz�`ֱ.u|���DuaP���pYѪvOR`�M�3*P�Q1Tl �oR�V�`�`A��B�N�m �>�b671TOC�a�QT!k�OPZ2���}���30e3OYߠREM��Rm�9�Oѐ$�reT�R�e��h�Fq/4�e$PWR�IM̃��rR_C�#tVI1S`sb�UD�#fs�SVW�B��b n�� $H.56�_AWDDR�H�QGr2�'� �
�R��~�o H� S��Q�4�_���_���_���SEؾA�HS��MN~�Ap T�0��_����OL����v���ּPACROx���aS�ND_C�����qٔZ�ROUP$���_X���@��1��25���?�4 ?� <@���?���?���2�AC�IO��W�D�:���J���1Sq3 $� ;�_D� �P�M���PRM_.��^�HTTP_�H�Qar (�OBJ�E��"�/4$�L�E�c��s �s ���AB_��T�SS�S� �DBwGLV��KRLÙ�HITCOU�B�G��LOF�R�TEM�ī�xe�a7f��SSQ ��JQUE�RY_FLA����HW��aQatZ�̯�F�PUR�IO �h����u�у��~�� �IOLN2�u��
@C��$�SL�2$INP7UT_�1$��i�1P m�D�SL��Qav��gߢԝ�=�s�=��5_�IO�F_AuS�Bw%0$L:0'�:1�q��U`|p�aaTժ�_��pHY�p ���y1��UOP�Ex `��>������hᣐP�Ã�^�`����x�!UJ	�y � � NEΩwJOG�g��DI�S�3J7���J8���7!PI�a���7_LAB�a3�������APHI� Qt��9�D�@J7J��� �@_KEY�� �K�LMO�NQaz� $XR�����WATCH�_� �s98��ELDb.5yn�E{ ���aV�(���CTR`@s����%RLG��|���DSLG_SIZM�� &��@%��%FD0I $;�Q2#�P=/ " _�+��@��Щ R ��P��S��� ��ťV" ZIPDU��r��N��3R}J����@P�A��]�d0U��-�L6,DAUREA��/�h�^GH0��!��BO}O2~� C�҆ӐIT�Ü>@��R{EC�SCRN�����D����'�MARG�2Ҡ�����N�"$����S3���W����A��JGMG'MN3CH����FNd�J&�Kp'PRGn)UF�|(�p|(FWD|(H]L�)STP|*V|(�e0|(�|(RS�)H�+��C�t�#y���1P#'G9U籐$"'�r�0&���"G`)WpP�O�7�*��#M07F�OCwP(EX��TKUIn%I�  #�2 ,#C8#Cl p!�p�� v3@���p�N�s�ANA�҉b�pVA�I��CLEAR~�vDCS_HI\T��Bu��BO�HO�GS�I�G�HS�H(IGAN; ��Mm!��T٤f�@DE�(4LL\�LC���BU�PR`���pT4B$1EAM�����7��#A�����pW��Ρ4�WOS1zU2zU3zQr�_�AR`� �����΁�esԲs�ID%X�P�r��O�P���a�VST?�RiY���a �$E�fCkW��&f9f.�DG�S��V�� L ���_�#�|p��U����וE��֕ESc�_ � �� .�x����c �MC �� ���CLD�P?�J�TRQLI��[����i�dFLG ���`��srAD��w���LDutuORG��!21r��vyxu���t���cд� ����t"5�du� PT��`��bp�t�vRCLMC�t}��y����MI����� d�)�QRQ����DgSTBP��P [��h�AX�bi�k���EXCESy���>�)M��U��O��dPXQ>��V��Z�]�_AW�\��������`KB� \�����7$MB��LI�I�REQUIRE�c�MON�
�a�DEB�U��;�L�`MA� ڰ ᛐ����q�;�ND>S��0'��ړDC�2:sIN�7RSM������@N���F3��P�ST� � 4n}�LOC�VRI��v�UEX\�ANG�R�Y�;�ODAQA��K�$t�1RBMF ��]���Y�b0�eǥ�C�SUP�e��F�XS�IGG� � ����b�wÓc:6�d���%c�?���?�.���DAT)ACWk�E��E������N"R� t��MD��I�)���@��-���Hp��ᥴX�!���ANSW!��`Q�1��D��)|��� n��� ÀCU; aV� px���LOj"�����5�W�3�E���U�M�;�RR2>B��� (E�N�A�q d$CA�LIa��GvA��2�9�RIN� ��<$R��SW0���)��ABC��D_J2�SEu�Y���_J3:��
��1SP���Y�P���3�"��
Y�J�J�Z՞r��O!QIM��(�CS�KPz��1oC��Jq(�Q�ܺՠպհ׎e�_AZ�rV���E�LQU��OCMP0s�)����RT���G�1���5��P1��9�f�G�ZE�SMG00}��Օ`ER���Å�PA �S(���D�I�)�JG�`SC�L����VEL�aIqN�b@��_BL�@Y����Z�J���������-x�IN�ACcR���	"x��f`_u�!�<���<�b܂�F���x�DH��t;����iP$V����'A$d�b�ȏP`��qy�B��H �$BEL��||�_ACCE��� �����IRCi_����ppNT�Q��S$PS���bLXP� (s�	1<w@
PATH��_D��_3..���_wQ �� ��rb�CC ���_MG !$DD���`�FWE�~���������DE�P�PABN6ROTSPEE�{Q�`��{QDEFb���XP?$USE_��BC%P��C�0BCY��Z�q s�YNA�A�p}yм�}MOU�NGRR� O��Q�INC�m���h�x���i�ENCS���d�Y�&��f�# IN��RI.%���NT�����NT23_Ux��`�A#LOWL�AA~0��`�a&Da0@Y�C���`���C,��(&MOS�@�MO��ǀ�wPERCH[  ~#OV�� �' �Q�#F�d"&�F��
�gm �@w�A. 5L ADw��v�)%�d*_6�z&TRK���QAY I�3쁏1.�5�3n�p�����PMOM B�h��sp"�W����0�3azR��DUЋ�S_BCKLSH_C.!E��&� ��-�?D�JJ���CLALBP'"�q�0܀|E�CHK�`�US�RTYJ�N����T:Seqr}�_c�$_UM����IC�C����C(LMT�_Lwp� T̱WE]&P[P !U,�5A�+0gT8PC�!8H�`|��2�EC�p�bXT���CN_��N���V�SF���)Vg�a	'�|�Q(2
e�XCAT�NSH������eq�
A
&F�/F�Z� P�A�D�_P�E�3_ �`���6� �a�3�d�E�JG�p���cO OG|�W��TORQUY /Ւ#�9� ?��"��� r_W�5�4C��<tP��;u��;uIC{IQ{I��F��.qaҐxp�� VC��0b�Z��r�1�~���s��uJRaK�|�r�v�DB���M���M�_DL��:2GRVBt;���;����H_L��b �i�COSv��v�LN�p�������d�@��mq׊Ō�q�Z����&�MY�����T�H��6�THET0j%NK23��`��㶣�CBe�CB��C��AS���mt���󌘑e�SB��p�GTS��(C�m�=���cM��ԃ$DU��@C7����� ���Q�F�s�$NE��ؠI@���C)���T�AX������h�s�s�LPHv�_�9%_�S�ңŅ ңԅ_��������EV��V����VʪUV׫V�V�V�V�V�H��E�²P��?aٸ׫H�H�UH�H�H�O���O��ONɹ�OʪO�׫O�O�O�O
�O�F_�����Ņ��Ė�SPBALAgNCEQԃQLE͐H_X�SP�9��ņ9�ԆPFULC�=�d�L�d�ԅ&�1���UTO_�@�eTg1T2����2N�A ��?�Ԗ��1f�D�5���1TP0O����,p�INSEG��!R�EV�փ "!DIF�y5K�1�0��1�� OB&�lAE��72�p?�A$�LCHW3ARlAB�a�5?$MECH��%�X���FAX�1PJTp��z���З 
��q�%ROB� C�R(2��Rf���MSK_���� WP ��_WR���r0�?{41	b4 2`0�1#JD0���IN���MTCOM_�C�p��  �� 8�$NOR�E$#���t����� 4�0GRr��F�LA�$XYZ�_DA��nC DE�BU�� ��t��u 0�$uCOD[AG ���2���0�$BUFIND�X2 ��MOR#�� H-��0����FB �0�JD$���c�QVPTAA�+�2G6� �� $SIMU�L�` 13�3O�BJE;ТADJ�US�� AY_It�A	8D�OUT�`����0�_FI�=@T+p4 ��X�3p3�A�5DNrFRI(CXT8E�RO�` E3q[0��OPWO�p'�}, SYSBUq�( $SOP��A�U�3�PRUN,v��PAC�D��℟0_� NR�X�A�B��PP� IMAG�[A-�G�P�IM�Y"$IN,��!#RGOVRDM�� ��P   #`W�L_`��an%�B�PRB5P�X�`QMC_EDT/ �� PPNq�M�"<OQ@MY19NQ+ �M!SL;�'� x $OVSL��wSDI{DEX�S��&�SP1�"V3p�%N 1q�0378�"<��$_SETp'��� @�0K2��AAR)I�� 
^6_��j7��1v1�5� �P �<T���`ATU}S@$TRCI�8H%�3BTM�7�1	I��$4NQ�3� '�� D-�E��"�2z�Ev��1!0l@�1EXE�0�A�!B*B��4S3�Z0.��0UP���9A$Y�' XN�N�7�q�$�q�9_��PG��� $SUB�1��1�1~�3JMPWAI,`P	3�ELOP�����$RCVFA�IL_CH��AR -���Q�P�T�U��R_PL�3DB�TB�a�R�BWD�V��UM�`TIGp�( ��4`TNL(`TjRRm���`
p	1	XQ� E�S�T�R�A�DEFSP�� G� L-���P_�P��SUNI#�7�PbmAR1@&�3�_L�IP�1�Pw�&�����`�� "<0��)�T"N�U�KETb(p��r`P^R&� h� ?ARSIZE���h1��naS� OR�3?FORMAT��TTcCO� ja�EM���d�SUX�2#�aLIOR&� � $��P_SWqIu�C5�cLLB&���� $BA̙`1�ON9AKPAM��0=y��BAJ5����2r68v��_KGNOW8cNrA�U9A"ߐDx� �PDC�ryPAY�[�t���y��wZ�sL�1��U!�PLCL_$� ! �s,qv�t�b"�vF�yCRP1O�z�2�tES���w�R4��w�tBASeE$�J�"W�_J�q
K�mA��fBu�4�r�qN�AX4P�`�AL_ � $��Qh 1q�!��C[�D:�sEfr�J3������ T� PDCK�� ��T"CO_J3�������
�hr���� ����C_YQ�  � �� �D_1
�z2�tD���n�^�x��m�|TIA4��u5��6[�MOMS @��ȓ��ȓ��B�@�AD��억��PUB{R͔������e#��` I$PI�$�QM�=q �wk�B1�yk���������iqRM�q�!Ħ~A�Ħ�A
��9d5S/PEED�G�b� �E�T��T�EP-��C��Q+�Q�ESAM(�E�����Ep{� m�$��  k�~@Ƕ�P_�ֹm��k�v{��ŵ��,H��ǳIN̚�c�� 1���B�W�.�W�wˏGAMM��1���$GET9" �D�;�u
��LIBRtcA�RI��$HIb@!_=!�0k���Eh ��1A����LW��4� +��X��7���wP���CEUv�[ �0 �I_b�xu�� L�������ȓu��پ�� �$Ј W1���I�0R���D\��kAT��LE@f�=q�1M�7�ୄP_MSWFLTM��SCRsH7�����!ؐ�~B�dSV&��P� A �����#S�_SAqs$��eCNO;�C�1fB<����� K�����S�C���hrǥ��m�D� a����  ���в����U!�C��������s ��cMJ�� � F��YLi�K���^SJ�|v!6O�K����BK�- ��OW���9���M$P��p����Dc$�"��1~B�`M��T2?� � $-�$�$W� �%ANG "�q� ����!� �5P&��o����c��#��X`O"���Zpz�`�@� �y�OM��+�(�:�L�8^�p���CON@�euL;�_�B� |� ���ș@&��@&�����m'X&��.��� (�0!%���`X$$�Pma�PM0QU��� � 8#`Q�COU���QTH�YPHO/� HYSf�`ES-r� UE� ���S`O�d�   �$P�@�Ŋ2UN��0b`O��  � P�p45�E��C�R�ROGRA�1A22DO445IT�Ё1�F0INFO�� �%0g;�1A�!O�I�2� (�SLEQ���1��0k6E1yS�НD� 4#`�ENAB"20PTION�C�T̢/G�T�CGCFA� @b#`J$P��<2����RdH0OBG�b\�E9D�@  � �{�K�q�3��E)�N9U�G�HAUT�ECOPY�qI0�L���M��N�@�K��PWRUT �BNV@;OU�b$G92DT�L��PRGADJ���bbX_ �R�$`pV�pVWnXP@nX[�pV�`Pz�N���_CYC"!R�GNSE�$ ��L�GO���NYQ_/FREQ0�Wb��a�d23L�p�b�PnQ8Ób��5CRE���#f��IF��s3NA���%?d_G��ST�ATU' ��*7MA�IL��YsIN��$L�AST�a���TEL;EMA� �GFEASIA�� ��H �b�1���f;B����I�0���R=q�!� LR�rAB+A��Ex0�V�a7vW�Cy��1�1U8�I0�pd�lv?RMS_TRs�� @��sr7�z��aktB��R�/ 	�b 2� =�_+� �ve��w�r� �fe�8�c�G�DOUa3;�NHC�RPR	 @���2GRID�1+CB7ARS��TYC�R'OTO㐾�³�&0E_[d!�P��B�Ox>D� � �0��PORa3��[���S�RV_`)˄ÆDI�T^�������砪�4��5��6��7���8�ZQF��A�~#0$VALURs����d�qE0F�U��� E��u1��aa��=@AN�㉒qa�R�@a��TOTA�L��1��PW�SI|J���REGEN����#XxxI3e%!���� TR^s0���_S��^���CVnQ�D��B8rE�cN��!��42��@ÓV_Hk�DA8�~���S_Y
�r�fS��AR�2�� <RIG_SE��ch�Â�e_80��C�_v�`�ENHAN=C�!� p�qEqqb�ý�INT���� F.3MAS�K��ipOVR�#P � N��`a
�_�*6���M��B[��f8��S�LG����� \ ���eH ���S,q�dDE�U��*7�Ő�%��U!�T�Ej  � (�7��҆�J϶�"cIL_M!d��P㈠�TQ� �Ë1rpj�e5V��C��P_��op���M��V1��V1���2�2��3�3
��4�4���ᄠ��`�����s��IN��VIB� �İ����U2��2��3��3��4��4�ؾ���#"�� �����%��׌ՠՌ�;PLv`TOR� ���INb�����  �{p��MC_F� 	���L����B��ڐM�IB���#� �1 �)���KE�EP_HNADD"��!��<p��C�_`A�䂁��H ��O�!���P������G���REM���쑥�;��R�W�U[de��HP�WD  ��SSBMo���G�1��2�� H COLLABu��a������4ؑEb�0IT��¸0��� ,� F�Lbq$SYNT��M�C��d��UP_DLY��#2DELAJ �nb�Y� AD��P ��QSKIP�� 	Ļ�60ODD���t P_60_2�g0^  ����		Q�	��	%� �
2��
?��
L��
Y�z�
9�Q�J2R�P*��CX]pT�SY��X]P��Y�1��� RDC��b�� %��@ReCg�R4ae�8�"d��RGEr@sl�:�FLG�!Pa�sSW�I��SPC�3��QUM_Yt�2T�H2N&�# L �1� �EFv�@11�!� l��`���C��AT4� ET1��7s"k0o4j!�@�Y�j!<3\�HOME(�"�P<$2D"�J/\/�n/�/�/�/�'3D"Ҁ�/�/�/�/?!?�'4D"�D?V?h?z?�?�?
�'5D"��?�?�?�?(	OO�'6D"�>OPO�bOtO�O�O�'7D"ր�O�O�O�O__�'8D"�8_J_\_n_�_�_R�%S��1�9 �q�=#$��pR�E���ٷ��LbݖJcIIOq�jiI�P��Gb�POWE��� �4` wo < ה ���b$DSB��GNABqՔE C�) �eS232Peܓ ���U�P�I'CEUQrt�E3 ���PARITáՑO�PB��FLOW�TR`�c�3����CU+pM��UXT�n���U�ERFACttC�Uѐ�b;CH�q� t����1_p��$����SOM۠9�A�T>�.��UPD�A#�`	T+`҃*�� �x�s�!��FA������R�SPqpQ��� }!�X$USA ؆��Y�EXmpIOH6��pU�YE��b_��0��B�#q`�WRp��_��YD�����VFR�IEND���UF�RAMδ��TOO�LȆMYH����L�ENGTH_VT�E��I���[�$�SE�`��UFIN�V_�@�5aRGuI���ITI�b��XX�	�J�G2J�G1T�U�D�d�u���_Â#O_p�py�ၻ��n�C	�zŔ��C ���ʖ �G���zr2�� @  9�qC���d�wu��ys�F� ���p��wX #�E_M�pCT^�H��f��<u�6�	�G#WV�z��G���Dh LOCK�~�U� ������=$� 2���~��D ��1���2��2
�3��3���:�����V��V=�"�=�F�V��!Ѕ�/������p�xṿ�����Prƻ���������E�������!��AC��PRs�!�}�S����`�Ec	��a�# 0 5�ؠ�V���ؠ���	������
zM�S��� ح��R�qda��$RU�NN�`AX2q��A⸀L�+"��THI�Cx� w �u��F�ERENg���IF��x���I����V��G1&�*Ԅ�1ٲ[��I�_JFR�PR���
��RV_DA;TA�q� RD�Z[ 
�AL� �xՑ �b{�  2� �S�~�`�	� �$ zZ"GROU���!TOT����DS}P��JOGLIYsN�E_P�PrO���\7`��bvK�p_M#IR�.䎐MQ�O�APp��E<�o��t���SYSE�ib��PG��BRK���v$ wAXIa  �������Ҽ�A����H�OBSOC��T�N�����16�$SV�1�DE_OPNsS�FSPD_OVR�4 ����D� �OIR+��PN�P,�F��l,��OV�SFa���d�$�F}�ja2㒓8��ҁibLCHH\RECOV�n���WE�M����RO�Ns���_���� 9@�9�VER��n��OFS9�C�Я�WDE���A����Rh���TRBq6aY�E_�FDOh�MB_CiMkS B��BL��.�u��8�V摁��p���]�Gv��AM���i ������_M�� [r�ec T$C�A��D��HcBK�q�vIO��q,�a��PPA �L1\D��bDVC_DB<���q �b���ja�1���3���ATIO"i`jqcp�U�� �efCAB�����J� �������__p�v?SUBCPU�b�Sv��`_��p"�`'�}���b"�$HW�_C� Ip���'ɣA�x����$UNIT��� � ATTR�I���"�CYCL���NECA�Y�F�LTR_2_FI`#��h��f��LP$���_SCT��F�_�'F_�,E2�*FqS�a��"CHA���-7�1�Pr�2RSD�  �b�����a�`_T��PRO�MFpE%M	`_���Ts2��� s2���5DI�&��tRAILAC4���M��LO�����5��������+PR�S̑{�dA�C�p	��FUN9C!��RIN됫�0|�@�DEqRA�@��� �C7`�CW3ARB�	BLƑ�G��DA�K�!�H�HDA`��AX�C�ELD�p �@S���A�@S�TI��`U�ѓ�$�<�RIA�q�bAF
Q P=��S��U �8���3MOI� P�DF_ꀔ��qHpL�M�FAE�HRD]Y]�ORGEPH�0���|� P�UMULS�E���`'���0J�(�JC�X�S�FAN?_ALMLVBs_a�WRNfeHARD����v�䐟p�@2$?SHADOW��0Ѐ�a�b��_`+q�ї�_,���vAU�Rx4\r?TO_SBR��e����j� ��A	sMPINF���!t6Q�'sREG���aDG�BP��V�p.�l�FL4�%!���DAՀ_X�P�CM��NЍY�B�V  ��� ]���$N��$Z�� �Ҭ����o� �|�EGK�����qAR��#���2?��wP��AXE���ROB��RED���WD���_F���S�Y��!���h�Sr�W�RIE��v� STRP���`��7�E�!�����a��B�����@CD� OTO7q����ARY����.A����#�FI��9�$LINK�Q����y�_���6���8�XYZ�bB�7NP�OFF
 �7�J+��B��yB��0���0}@��FI� ��Є���yB
�_J ��5�����`Ȅҋ8��H�TB�b��C0x�DU �9.AETURa`XgSW����rX���FL�z���#�pu�Y���3x\��� 1��%K�M����31�DBp`%��`'2ORQ�6 �ѳC��}�DB��>��P���%�����\q:�OV	EA���M90=ѻs[� �s[��rZ��`X��aY� � X�O�~@91�P��B� F����=�S�B�_��0�s����ER�A�	EBE��� QC"�Aб�����E�2��Q&QAX���Q�  �!�|�A��+a��� ��@@��O���n������N���1����`�� `��`��`��`�� `��`��`��`��!��� �Rg�DEBU�#$�A�c�2��3�ABGE�;�9V�" 
�Ҷ ���z!$�
�$��$� @A$�O�$�n�$��$��N��T#��R����LA�B���� �GR�O0��l� B_ �1	ƞ�>��`���p����a	�ANDà�E ��<���aF�  ��q��Z�Qi�� ;�#NTq`�cR�C�1=��
��	 �pE�RVE���p� $�q��@A�a!��PO�`X �����Q��p�  $.��TRQm�
��Q�2����R2�oP~@_ � l=����fERRҒ�I�V����gTOQ����L%��Ď�z�0G��%%�"��?�!P � ,��2 �뺱RA� 2� d�D�p� 7 �p$O��2��PvµOCQ� ��  YCOU�NT���FZN_wCFG��� 4� ^v2T�d�"���m �W k!
E�s� ��M�08b�����X��0�FA~P���V�XA������0����O A�P�b�pH�ELkpN�� 5ސB_BASN�#RSR]vm@;��S�!YQB 1�B 2�e*3e*4e*5e*6�e*7e*8�5!ROaOGP� �:�NL�q�)�AB��@C AC-K�INT80�s�U�``x1�)_PUXA��b�2OU��P�@�^x"#�y0��b�TPFWD_KARlLfpZRE���PP��&Q�@QUE]zRO B�2����`�aIb`��"#8�$C0Bv8�SE�Mա�6�`A�S�TY4SO�0�dD�I1�@r�1aǿQ_�TM�sMANRQ�AF8�END�d$�KEYSWITCaHS3h1#A�4HE2��BEATM�cPE��pLEks1���HU�g3F�4h2S(DDO/_HOM�PO�a� EF"�PR���rS�����v�@OaX �O�V_M���`pPIOcCM$��7��v##HK�q� D5�$_w�U�b�2M�p�4�4�%�FORCcsWcAR�R�p!%OM�p � @��˓�`UU��P�1�V2�V�3�V4��O�x0L�R��^xUN�LO.0�ddED��a  �$$C�LASS `����.a�p�P7`#`Sܘ0+h�P��?aIRT?�,o>`�AAVM��K 2� je �0  �5�5a�o�h�o�m �l	�m�pk`!��o2v7u�lV}�b�ah���t{`B�S4�� 1Li�? <�� � �2�D�V�h�z��� ����ԏ���
�� .�@�R�d�v������� ��П�����*�<� N�`�r���������̯ ޯ���&�8�J�\� n���������ȿڿ�h����rC`�AX��� `���s  ��%�IN.�@�$�PR��0XEQ�}�`�_�UPMIl�ja{`L�PR ji`��tLMDG �g��`��PIF 	�k`d��0�B� T�b�߅ߗߩ߻���, 
���n��o �0�B�T�g�x���������yNGTOL�  �{�pA  � ��
�{`Pd�O �� ��=�O�a�s�6b� ��u��� 2b������������&@J4Z������ �����*�<N`r��zPP�LICA�1 ?�je}�����Handling�Tool � �
V8.30P/�58��
88g340��F0!�755����7DC3����None�F{RA� 6*-�  !�� TIV(qŵ>��#UPn1�R:b\�PAPGAP�ONf`�.za� OUPLED 1�i� /03?E?W?��_CUREQ 1M�k  P�a7a<��n�?�d}��33b{9b ��Ƨ4H�522�:HTTHKY�?Kx�? �?ZO�?6OHOfOlO~O �O�O�O�O�O�O�OV_  _2_D_b_h_z_�_�_ �_�_�_�_�_Roo.o @o^odovo�o�o�o�o �o�o�oN*<Z `r������ �J��&�8�V�\�n� ��������ȏڏ�F� �"�4�R�X�j�|��� ����ğ֟�B��� 0�N�T�f�x������� ��ү�>���,�J� P�b�t���������ο �:���(�F�L�^� pςϔϦϸ�����6�  ��$�B�H�Z�l�~�0�ߢ��6s5TO��/��#DO_CLEA�N�/�$6�NM  �� a?��������g>DSPDgRYR=�p5HI� `�@q�8�J�\�n��� ��������������m8MAX�����17.X�-!*2-!�"PLUGG0�*3��%PRC��B^�"b�'��O���^
�SEGF� K� ��^�p�8J\n8���LAP�( �3���
//./@/�R/d/v/�/�/�/�#T�OTALPy	�#U�SENU"; ��8?�2s0RGDI_SPMMC� o1�C�@@@
�"4O��5 3_STRING 1	�+�
�M� S��*
�1_ITE;M1�6  n�-�? �?�?�?�?OO'O9O KO]OoO�O�O�O�O�O��O�O�OI/O SIGNAL�5�Tryout� Mode�5I�np?PSimul�ated�1Ou�tQ\OVER�R� = 100��2In cyc�lEU�1Prog� Abor[S�1~;TStatus�3�	Heartbe�at�7MH F�aul�W�SAler�Y_ oo$o6oHo�Zolo~o�o�o  �;�?�o�o );M_q��� ������%�7��oWOR� �;o��o I�������͏ߏ�� �'�9�K�]�o�����य़��ɟ۟�PO �;�Q�����6�H�Z� l�~�������Ưد� ��� �2�D�V�h�z����DEV���*� ��޿���&�8�J� \�nπϒϤ϶�����������"�4�PALT�m[ч�5߃ߕ� �߹���������%� 7�I�[�m�������I�GRI3 �;�� s���'�9�K�]�o��� ���������������#5GYk��� R �m��}��� %7I[m� ������/�PREG_�H �!/ o/�/�/�/�/�/�/�/ �/?#?5?G?Y?k?}?��?�?�?]�$AR�G_o�D ?	�����1��  	$�V	[
H]
G��W+I�0SBN_C�ONFIG 
��;IQHRCACI�I_SAVE  �ThA_B�0TC�ELLSETUP� �:%  O�ME_IO]\%?MOV_H�@�O��OREP�_�:U�TOBACK�A�SMFRA:\5+ _5&�@�'`�P5'dX�= q^ ,H5-��_�_�_�_�_*o]T���0oXojo|o�o�o �o5%Eo�o�o& 8�o\n���� �S���"�4�F� �j�|�������ď֏���ۏ ��$�6��H�Z�!_INI^���U[E-SMESS�AGw@���A�0��ODE_D�@zFDV���O��ǟ-SPAUS�'� !��; ((O�2�1��Q� ?�u�c����������� ����;�I����?TSK  
�d_<j�0PUPDT�����d��ԖXWZD�_ENB��WJ��S�TA���1���1WS�M_CFO@�5�]E�7�GRP �2� 	BB��  A���9XIS>I@UNT 2j��C � 	z���A ���Ϭ�����	���-�p�=�c�f�MET� 2u�PNߧ�J����^�SCRD�1J��P�EB�� $�6�H�Z�l�~�]_5*Q{I��������� (���L���p������������1�k��73QGR�n����	UP_N5A�@�;	3T�_ED��1�
� �%-BCKEDT-���J��&U /dD�@-3Sz
5*,B&o�Fs&/  ��2�K �wʹ�E��	�-3�X5/| �/|/��k/�4�/$/?H/��/H? �/�/7?�/5�?�/ �??��?O[?m?O�?6LO�?�O�?��uO�O'O9O�O]O7 _�Oe_�O�A_�_�O_�_)_8�_�1o��oxo�_�_go��_9�o o�oDo ��oD�o�o3�oCRS_���]���Ug��	 V N�O_DEL'GE_UNUSE�%IGALLOW� 19	��(�*SYSTEM�*��	$SER�V*¯�Ȁ�REG�х$��ȀNU�M���	�PMU|t���LAY�����PMPA�L��J�CYC10�U�h�R�V���UL�SUH�
�j��Ӄ�L��ݔBOXOR=I��CUR_ʐ	��PMCNVD��ʐ10~�0�T4�DLIȰß�ˋG$MRߎ�&�&� ϲ����̯ޯ���y�	 LAL_OUT� k��(WD_ABORo����m�ITR_RTN򩷀��m�NONS�TOM �� ԸCE_RIA_I�������˰F���U�c���_L�IM߂2` �  N��Nϯ��<��m�`���� A?Ϡϲ��ϯ�
�����p��PARAM�GP 1U���Ύ�O�a�s�2�CO>  CV���f��Qz�ߵߗЇ�Б��U��Р�Ъ�д����٢���������C����ǀ Cї���+���?�ɲHEC�ONFI�w�E�G_P�1U� 49��������������E�KPA�US�19� ,�uG�Y�C�}�g� ���������������1U?e�!�M~��NFO 1(�;� �=������� D��B��D�  6������ ˰O����ǩ�CO�LLECT_�2(��pEN`����\�INDEx�(���!�12�34567890���������H,��)'/L/�|&/8/ �/�{j/|/�/�/�/�/ ?�/�/?e?0?B?T? �?x?�?�?�?�?�?�? =OOO,O�OPObOtO��O�O�"� � �ɶIO "�����O_a_s_l�_WTR�2#]�(�8Y
�O�^P��$,]�Z��Y_MO5R"�%� �9�Fe �Fi^oLo�opo�o�k�b�#�&-mB�? >�>����a�Kt��A�PM(���a�-=�Oas�� ������^@
�����` *]c�PDBO*����Ecpmidbag�C���U�:�Ձ�i)�p/���S� G ��,�l�-�,̏����9��v�������1��gX�^�)� 7��fM��w���@ud1�:˟���Z�DEFg )o7S)ߑ�c�buf.tx�t��M� �p_L64FIX +� Q���˓�د��ɯ ��2�D�#�h�z�Y� ������Կ�ſ
���.�f�x�_E ,� �l�~ϐϢϴϬ��p�IM�C-�]���6��>���=�L����MC&c.D�SdF�'�%d/5�!�`t���B!!� ����߲�����n��gM1�\D�y**��~**�}���`U�x*��C�ÇЯ��BDw�4�  E	3��Ee��3Ec��Et�� F�3E޿ŚF�B���F����F�YfF��% G�� G	ڳH�3�?�  >�33� ;���a�v  �nf��q@35و���b�pA�a�<#�eDQ��7���F��RSMOFST c'�f�G�T1#`uDZ�2!���Q,�*;�0�R�L��?���<�M^��TEST�0���FRz3SMx�C��A��*e�h��| C��B��3C�pn���*�:d�b2Iy4�<2T_�PR/OG ,k%^��/%PNUSER � �1��KE�Y_TBL  �-e1]�(��	
��� !"#$�%&'()*+,�-./�:;<=�>?@ABC�G�HIJKLMNO�PQRSTUVW�XYZ[\]^_�`abcdefg�hijklmno�pqrstuvw�xyz{|}~�������������������������������������������������������������������������������͓���������������������������������耇�����������������������A� LC�K#D#STA�Ti/0_AUTO�_DOG㺒�+IN�DT_ENB�/ a�"��/�&T2�/�6STOP�/�"S;XC� 25K�p�8
SONY �XC-56Q{�}�p�@��͞b} �PАX5HR50��-tx?�>|���?�Aff�:�O"O �?GOYO4O }O�OjO�O�O�O�O�O��O_1__U_g_�\T{RL� LETE6� �)T_SCR�EEN -jOkcs��PU0�MMENU 16� <O\�o ���_oIo��&oLo�o \ono�o�o�o�o�o�o  9"oFX� |�����#�� �Y�0�B�h���x��� ׏���������U� ,�>���b�t������� П	����?��(�u� L�^����������ʯ ܯ)� ��8�q�H�Z� ��~���ݿ��ƿ�%� ���[�2�Dϑ�h�zπ���ϰ����b��S_?MANUAL"?�Q�DBCO� RIG��Ws)DBG_ER�RL� 7�[������ߴ��� O�NOUMLI I����dD
O�PXWO_RK 18����&�8�J�\�n�DBwTB_�Q 9<�����K,�D�B_AWAYW�^��GCP D=����_AL �/��SҡY!0�UD H�_q� +1:����0,R0�`T���A�~���_M� �IS� ��@� ��OoNTIM�W�D�����
2#�M?OTNEND'"��RECORD 1�@� �����G�O�N<����z ���G��N r'9K���� ������#/ �G/�k/}/�/�// �/4/�/X/??1?C? �/g?�/�?�/�?�?�? �?T?	Ox?O�?QOcO uO�O�?�OO�O>O�O __)_�OM_8_F_�_�NIO�_�_�_<_��_�_�_'o�N��� (o_oqo�_�o�o�o�o�N\���o�o=p�oH�o��B��p ��(�����N%��K�]�����TOLERENC���B����L���O�CSS_CNS�TCY 2A~� h���Џޏ�� ��&�8�J�`�n��� ������ȟڟ�����"���DEVICEw 2B~� �� r���������ϯ�����)�����HND�GD C~�C�z<���LS 2D\�;�����Ͽ�����=���PARAM E/��i�����SLAVE �F~�J�_CFG� G/�)�d�MC:\��L%0?4d.CSV(��c����A ��C	H��n�n�)��=�
[��)�-�Z�j�X�<W��JPъ�C��_CRC_OUT H��<�+ϑ�?SGN I���
�05-MA�R-25 16:�01����て Ze�7-�)�)��*঴\�o���Im��P�uG��=��VERSI�ON ��V3.5.20���EFLOGIC {1J% 	���* ������PR?OG_ENB��\��ULS�� ,�P��_ACCLI�M����Ö~7�WRSTJN��0��)��MO�
���x�INIT �K%
��) v�O;PTp� ?	�����
 	R57Y5)���74��6���7��5��12����6����TO C ��@���V��DEXd�do�x�~�PATH ��o�A\����IAG_GRP �2PI�|O�	� E7� E?�h D�� C�� C ��B���C��nk�p��C���Cm�B�N��BzoOB�)��Bk�f�383 6789?012345����B�  A���A���A��A�O�A���A{+As��Aj�RAb?JAY% x�@���p��G!���A�p�p��B4�h���x�
"�����"�Q�A����A���A����A�� ��h�Ax~�Ao�7�Af9X��?$>��mF/X/��h����(�"_�AY��;AS�TAM��^AGdZA@��A:bA3�%A+�-A$����)�/�/��?�*@��;d�6���@�{�@u�-@�o�@i�7@�cC�@\�j@�V{N?\0�5?�b?t?�??@_���@Z^5@T���@O�@IG��@C33@<���@6�+@/<@(�`J?\?�?�?O�8�s� nE�@h�@b�!@\�0�Vff@Pt@Ih�s@B��@;�bOtO�O�O�O�'6] ^_p_N_�_�_0_z_�_ �_�_�_$o�_�_
olo ~o\o�o�o>o�o��C�"�!30�2KA�@^>�8Q�r��R?��  *u^7����Fr'Ŭ5AFyRu^@�p�nvF�@@�pppE�@[ �Ah���uC=+�<��
=T���=�O�=���=�<����<�p�q�xG� ��?� �C� � <(�US� �4jr�D@����,"�A@w�?f�o X��mf���������� ԏn��
��.�@��i�?#�
b��\�>�pn�^��G���G�^x���R����^8 Pۑ�5甮��CnB�AL]_u��&�P;�'f�d��aQ{����dD�  D�  C΍��̯ޯ 8����VʠǯD�ïh���� ��3+��Q�ҿ����� �,��P�;�%ZN�D����CT_CON�FIG Q-|��#�eg��� STBF_TTSd�
����C�V�:���MAU^��~��MSW_CF���R-  _ ��OCoVIEW�SY�i�����߽����� ���G��.�@�R�d� v����������� ���*�<�N�`�r��� ��%��������� ��8J\n��! �����"� FXj|��/�����//j�RCR�T�e&�!�,.V/ �/z/�/�/�/�/�/��SBL_FAUL�T UI*n�1G�PMSK��$7��TDIAG V���e�2�UD1�: 678901�2345�2��?�P �Ͻ?�?�?�?OO)O ;OMO_OqO�O�O�O�O8�O�O�x �>�;��
�?%_��TREC	PZ?l:
z4l_?��? �_�_�_�_�_�_oo 0oBoTofoxo�o�o�o��o�o�O_/_UM�P_OPTION�>*qTRR���!9�KuPME��>Y�_TEMP  ?È�3B�Пps�A�p�tUNI7���şqF�YN_BR�K WY�)8EMGDI_STA�u�&��q�uNC�s1XY� ��o7�*�~y���d ������Ǐ ُ����!�3�E�W� i�{�������ß՟� ���r�,�>�P�b��� �f�������¯ԯ� ��
��.�@�R�d�v� ��������п����� �%�7�I�[�u�ϑ� �ϵ����������!� 3�E�W�i�{ߍߟ߱� ����������/�A� S�m�w������� ������+�=�O�a� s��������������� ���'9Ke�[� ������� #5GYk}�� ����/1/ C/�oy/�/�/�/�/ �/�/�/	??-???Q? c?u?�?�?�?�?�?�? �/O)O;OMOg/qO �O�O�O�O�O�O�O_ _%_7_I_[_m__�_ �_�_�_�_�_Oo!o 3oEo_Oio{o�o�o�o �o�o�o�o/A Sew����� ��_��+�=�WoI� s���������͏ߏ� ��'�9�K�]�o��� ������ɟ۟��� #�5�O�a�k�}����� ��ůׯ�����1� C�U�g�y��������� ӿ���	��-�?�Y� c�uχϙϫϽ����� ����)�;�M�_�q� �ߕߧ߹���E���� �%�7�Q�[�m��� ������������!� 3�E�W�i�{������� ��������/I� Sew����� ��+=Oa s�������� //'/A7/]/o/�/ �/�/�/�/�/�/�/? #?5?G?Y?k?}?�?�? �?�?���?OO�? K/UOgOyO�O�O�O�O �O�O�O	__-_?_Q_ c_u_�_�_�_�_�?�? �_oo)oCOMo_oqo �o�o�o�o�o�o�o %7I[m� ����_���!� ;oE�W�i�{������� ÏՏ�����/�A� S�e�w���������� �����3�%�O�a� s���������ͯ߯� ��'�9�K�]�o��� ������џÿ���� +�=�G�Y�k�}Ϗϡ� ������������1� C�U�g�yߋߝ߯�ɿ ۿ����	��5�?�Q� c�u��������� ����)�;�M�_�q� ������!������� -�7I[m� ������! 3EWi{��� �����/%//A/ S/e/w/�/�/�/�/�/ �/�/??+?=?O?a? s?�?�?�?��?�?�? O/O9OKO]OoO�O �O�O�O�O�O�O�O_ #_5_G_Y_k_}_�_�_ �?�?�_�_�_�_'O1o CoUogoyo�o�o�o�o �o�o�o	-?Q cu���_�_�� ��o)�;�M�_�q� ��������ˏݏ�� �%�7�I�[�m���� ���ǟٟ����!� 3�E�W�i�{������� ïկ�����/�A� S�e�w���������ѿ �����+�=�O�a� sυϗϩϻ������� ��'�9�K�]�o߁� �߭����������� #�5�G�Y�k�}��� ������������1� C�U�g�y����߷��� �������-?Q cu������ �);M_q ���������	 /%/7/I/[/m//�/ �/�/�/�/�/�/?!? 3?E?W?i?{?�?��? �?�?�?/OO/OAO SOeOwO�O�O�O�O�O �O�O__+_=_O_a_ s_�_�?�_�_�_�_�? �_o'o9oKo]ooo�o �o�o�o�o�o�o�o�#5GYk}�_ ��$ENETMO�DE 1Y�U�  �P��P�U��{�pR�ROR_PROG %�z%�V�&���uTABLE  �{oe�w�������rSEV_NUM� �r  ���q���q_AUT�O_ENB  ��u�s�t_NO΁ �Z�{�q�� W *������	��Ā+�*�<�N��HIS���Q�p�_ALM 1[�{� ��T��P+O�˟ݟ���%�rS�_����  �{���rj��pTCP_VER !�z�!�5�$EXTL�OG_REQk�9�ቼ�SIZů���STK����~��TOL  �Q{Dzs��A ��_BWDJ��؆K��ԧ_DI9� \�U��t�Q�rU�STEPa�s��p���OP_DO��qF�ACTORY_T�UNk�d̹DR_?GRP 1]�yށ�d 	e�#��p��x����� �n��So �k� ���W��i�z�d� �ψ��Ϭ�����	�����?�*�c�N�@����@�!�?Ơ�s@+a�j�
 E���R��j��x�d����E7� E??p D����L��D�%��  Cμ��K�B�  ;��  A@E�o�@U�UUc�UUo�&�>�]�>П������E�F@ F�5U��{�L����M��Jk��K�v�H�,_�Hk�{�?�м�Q�9tQv+�8���6h�%7��{�T���FEATU�RE ^�UK���qHand�lingTool� �� rodu�Chinese� Diction�ary��LOAD4D St���ard��  ND�IFAnal�og I/O�� � d - ��gle Shift���F OR��uto� Softwar�e Update�   J70 m�atic Bacwkup��art �Hground �Edit���70�8\��ameraz��F��D pr��nrRndImMޤ�PCVL��om�mon cali�b UI q.�pc�nf� Mo�nitor��ws�et�tr��ReOliab	 ��jp �Data Acquis������ Diagnos�D����� Doc�ument Vi�ewe���
P�C ual Ch�eck Safe�ty� act.�Enhanc�ed UsGFr�w ��\weqpxt. DIO � �fi+ t\j7�endxErr� L*  � �{'s  ��r��� :���T "� F�CTN Menur`v���t I��TP In�fa}c%  48\� �G_ p Mask/ Exctg�� �o��T Proxoy SvH  5�p��igh-Sp�exSki� "� #1��#�mm�unicC onsn�apd�!ur ������"con�nect 2Pd�in� ncr sgtru�� I �KAREL Cmod. LE uaG"�t\ia�%Runw-Ti�Env�z�"K�el +G �sE S/W�?Licen��[�GER  �Bo�ok(Syste�m)�� R5� M�ACROs,x"/gOff� �Pa� �MH�- �: \ac�1MR� �)���MechStop�V!t�  ��0i8���Mixx��dE ��
� �0od
 �witch��Lo�a� �4.�6 k� G�1�3OptmpUHM GGW filG҅ HF��g�' p�mfO Multic-T= i�4pa�PCM fun�'�{3M"Po[�D zQV�HRegit0}r�   mpo� �Pri@F�K _�fcs W g Num Sel�5��� |DS� Adju� P���`W
 4 S|XtatuQ/bUC��� RDM �Robot��sc�ove�� cctNO Rem�0�n��<�SServH10@�#CTXPSN�PX b<2�� "�K9$`Libr����564@e�� X�4H`ZUSoY0t �ssag�E�~� �"�1�VVLO�b/}I- pc
�`�MILIB�mchy1o Firm+p�8� �b"Acc` <hXcTPTX�;��<� s Teln�0�m�}B��5��4Tor�qu
 imula��}�Tou7@P)a51��m�T_ ��QC&V ev. o�cleUSBg poU � iP��a@WdUSR E�VxP+Unexceptx�P�D{D,{f}VC�r�"�"�2�sVD��j�cV��Hk uifoV�S?P CSUI�k���XC�6X`We�b Pl�V��9pjxăa�+64.f���^ r>�T�v�
J�57À�vGrid��Qplay 76� (��`L&iR�;�.��K�\0ARyC; 4 120i��>L#AsciiV!eRpDAG�d��UplE@x��� �@CollW�;Gu�� of^QޝPI   1�s� ���t�0t8FK���Cyr�p  2*Porie�  ld�aFRL��1am͉ RIN�T��MI DevfO0 (&ax2 ,�0��A/�rb�@as�swo��9��64MB DRAM�
�IO" ��FROnƫ
! ��rciP'vis���qG`���Welds cia�l�40BW��el�l��a�BW�sh�/���"PH�cXEw'mrwH�( p�v{��ty	 sPR�"wm0�t!1m@.]��P ��P��'�8�D� %2b a���r �P+��r�Pb� q�drT�1� e�COL��S�up�r�ARged� OPT "W�8s�H��; cro�V C! � �SHe[�  � 
gq� �uestY  ��SS��e��tex;`LO S�p$![��E��bP�@ �4Y|CVirt�W�S��PPdpn��x�e~��e���y\ߕ�jui.x����ߖ� аߕ��51 J����(F9r�ߕ�II)�ߓ�on��!���M!=�ӈ	QY���f>�t���mfV��լ���Ҍr�� ��?���&P�3����Ҭb9���eie�߽�n\p���\R���ҭ`A��2�p����O!
!����O��j�7 J5�����5�ӝ1Q��\ar�7���XPR���k "��}��b����`9P���lnko����`1��RMJ�����;���M�����H5�4���883]D#ER�N��Ffh�FM/el���չ1d/ ������d0�/��|B �/�( �/��<��/��9p����.fd�/���ASTC?��616<�/��g HS|?z��as����j����?��0�?c�r AW$O��!`��%rzP]O��t\a[�U5�` �O�$�a�O�ҵ��O�0���O��.EN _�D8�`<_��ite_?���v t_�� aO��IF{?�Ԉ`����) "s_�Epa��O-�>n1!Ot.IvTo5!�_��F���o^837�o*QogW-���o�/��X@�PDT4��_�ԓze�OHf4�_\7	9���MN������f�tro9?6�x�9i0���J59L��%����Ak��P����_p�o�Fp_-o0�@�?(�f1'?�pm_d��O���ٟ�O.�pe����m\�A��/_���j�'2.p�͆cW_��֮͠c�a/\ Ry8���(Las$����O_���0x���bo��<����-�̿"%� ���K��/?�siaf<Ϟd�?�NT+���Se����//`�C/�����'37��fiUf\����$SG���Ԁ6���RDYaLS߱�oI�omw��_#�ps0����d�hVmj��93����E�ogW�P���ch\?�I��ퟓ� 8�o����rvi7�]�S�/������V(st�,��F���@�tl��u&5/����Td
�hWi��ݶSe��6O��sr��	��! ��y8P`��dr׏�o3PRI����a�O�/	X/��spr�ߕ��擇Li?/��3 H�6x/�d94'��6�3�q54 H�/v6353�/r4 H���&0�/�'��� X?v�72�Ie?�g13$;?��7�/58r?�'�6�/��Lo�_��t �ͅA�ϐOc�m�osK�!����O�����,�O9��O�OS�ua�lP_��8�?a_�^@gs��_��wr+��j83�?!�_]�&��NDSO-�f7O=��!�Y�ad�O9k1l�o�s_#1�o���ip#�-Et�op�RI�N,��/I���V�A�=SE_��0�
S���Z 0+ͅcmg�Z��0 4@�"�ut[/�of��`�M�r����@�����596O_��4DЏ��U��#o(� I�c5%r_����e`���G�������c���AL"���lga33_U�oy� -<�t
��	e�@t���RTU���h�z�xo��vo;��'O�52 ����4��'�2Yu\�� vOA���42I`FĿ
d -�ݕE��� (o�[��"E3�yo��Wel�_��������WMG��Ϣ3aP@�Ϣ3wm�g[����߂�- ����On�45�?�fCqMk�IO��  �� �������1���2�g��y� R�;�Co���4(S�`�⯔��Ġ��3IF���� 1!(�z�0at��cNT��q���R8��8i5�l82\��� O��W?��˿ݿ`￘��7��4SiZ/`<��=�K�!�cl��i5\sw/�S�AD̓��CVt�Dt.�Q�mt�_�e����V�-V�  /6��Nlo��1��\�O�/�C �/�4 �/�i`�e/�/1_��62˟2��o�/�eJ7���erv�?�) "�?�svh�?
o�N�� �?�.p[�tvshmoO�U749LO�R`r��Outl$O?�t\�?��j�_��//�/h_ mpcL��y�9\KO�j�_0�/�_�uXP�/D�cH8gO}�oOnn�O�%N�߬u�'o���np]`���oRCM�o�un�_��$./�_#��m  �H552�a�be�q38BSGR78�p�q�r0���libJ61�4�cATUP��@rmc�p545�zPsgt�r6��VCAM�3wCRI�p\rc�p�CUIF�  �q2ީptd.f�NR�EN rco�p631  - Pr�p�SCHV� Di�DOCV>aIF�L�CSUJ18�0��p1}�EIO�C  ��4�p54R�pR�`4�9�pgm�wSETf�Sta�q^�qlay,�p7�q��0MASK~�SPRXYZa�ap�7f�C�pH'OCOC��3.3�r6�p\c΂51�p���qapp.�q39�f�j50�q�us�t3�LCH��A`
?OPLG�1"��E�� "L3�MH�CR  08 (�ĀS@�Reg��C�S�p�1H��p��q5��p08\�pMDS�W  URGw�MYD���sOP��\!�MPR�ra�4�Հp!�o�f��p! p���PCM�H��R0БPath���p@aDH�ՀRm����pTP�ܠ�Հ816�50��pg��āS��ol�,�9Ղ:�FRD��p(Q�pMCN��c�c�H93�pLN=P��SNBA@�r�SHLB��֑SMnx�lrn?�63�p���q2�pL�HTC<�pX�TMILVs�r��T��PAu�Y�s�ȡTX>aEN��E-LU�th��0�@`�8�qHѰr9��`ρC95�p �Հ7���UEV��adin�(�C�����pUFRvI�eeO�VCC�p�t�VCOY���VI�P��spd�[�I�^�p�X͡tsπW�EB�p��?�HTTv�p L2�R62�p7Coo?�CG��d��IGt�
PR�I��PGSN ng��IRC��ne n��H84�prd6��R7��@�R��L�5�3�p\lcl�q8^�pD" #4�6M�� ��52�8�R6�59��|�5�r dK�R649����r89�YpS�D06�p1�zk�Fc�VG M�v��, ��AWS�p���ðCLI�J6�43H��p����u�z�dҡ���pGD��ScTY��$��TO������q6�<q|� �g���<�RSY�-@��R�68�p�OLp�3ι�OPIɰģSE[ND�guG�LP��ݠ�pS��T�ETSɰy�c��2!§�-��U��FVRu�43k !ıN��ry:��ytonF�yt Lo�a��D (S��di��I�0�֙���p��ytt\sg��g ="�ր6���L�yt\str�ոA��<�@��hk_t���yt����es�լr��{j7��mon.��(�A��d@6��s-@����yt46\�`Q��b�qh3��zDll���<�&Dc�`�$rt {������yt��w��x�U�Ӑh8��nde��AxV絰�����N��ͰH��epe!n���yt�T��Ģ���ob3攢��h8�9����p��Pv�e�d~���4 J7R805��0l��ձ`"t644�����G II���r�p����"S��#л%��w594G�tom��:�!�R J���l ��Se3�ar3�E�t32�%�QsysG�F ���������etr��urn�k����20�x718���'�rn6��l���\jtET�v�
jo��ta.C��gr������� 0���<���ge���017��2�yt�yt75b���k'���]7 "P��T`dc��) ��	�`���r��1%at�b@O���p��daW(?�4tv/ 4oh��c�8}���s?yR�?�=l�ogm�?�;ild�?1<d�?N�@���H0@O�M���p1|O��;x@���ytV��1����O_�	8�aicC 2�9����C��7��6�E �� `E?k3edg?y=wm�`O�Rhl$_�2G&heh>�m_��7�5l�O2 24O Oaw4OJmsdh\o�;dh2����osqz�o�kl@���o�o��:��+F�cet�'-�6J8"W<Q��1 (F���pbDa�0��fr{F�� �� �f22.fv�FusS�pkg�M!INgD�x����,��u��o�{��5s22�xsiRC��n VM��^�99�2�W� ��J9�b��st�'T��O 92\�6CMR/d#Z��O;��ݎv'���t�mF����f8�va%t��t+9>e��6ft"/��z_v(��ɟ?�4o
���,���կK����vs�w�8��Dni�o��lb��蟮���p��W�\���vsmTڴaz�"����οD��of���ow�L(ώ�slw���f����e�w�����*�vrh�ys�+N3GeN��v�Y25:�oad��(Na�NJ?��nd�� "NwV � ���@s����rrd�6`��le&���C�U�4;��Ok7\��8���1rk&,��gl��P�b��g�Gt��il��������  e P2^���38��r ����0~��J614�?ATUPj���545����6F��VCAM���CRI!7� , U�IFB���2��an=s��CNRE�'��631��RI��S�CH�u65D�OCVN�ns� C#SU�T|���0��HA�EIOC% �"��54��R69�65\� ESEAT�W�����7� Cu� MASK��t 1PRKXYUJ N 7��n��OCO�om�513r�,,�����<� ��98\t����,]�[39�v!���oftwLC�H!g�OPLGZ:�950ai�P�]P��e f,S2�r��CS�􈑼�g_lo��5r� �pDSW6��r70<!Pl D�KOPP4�PR�QS01� n Adp����X#PCMA	a ��0�%����vdv; �A
CTX��0��1AGDIG� �!H z,S�r723��q9AU�+ FRD!�h#RMCNr	H9�3��R2SNBAz"�C+ SHLB�	CSMp5�n m�wJ52�HTC��ިTMIL6�Seh���PO�0PA�{86*TPTX�V�R�0ELA4oolQ,��� P��8���\sv���qSR�VT��95Q$9�5A\et� UEV�@a\AC!]�[AKFR!r��C!wol.�VCO�\�P��VIP�4e�ڟ I�t34[SX|���WEB���@(�1T��,�l2�tQ, G�Eg\t�kIG�E#@`PP�GS"�PRC�4"7TAN��84��#[R7�taQR�(�
R53�tRJs68��R66av52a- E���R65qr Im��5a��l4q5�73��U�D06D�5`M,0�V�E6����WS!  m , LIQ40�A��Pf9MS�S�ni�@^`���SST�Y�4597[TO^��76 J��6�5�x��P9 (k O�RS�fer@R�68��C���\sun["I1TCSN� �S� 6׼�L�Ecs�n.\0�f �bET�S1TX�2E���0C�Pah#FVR�E6�6 IPN�5���|yCa
@}xBx}x��|yMG" |y<��|yg_cc|y"}xcmg_|y��yGvth|yR}x3(��,�>�P�b��z1��z!� cv|yon T�|yh"}xhr}x�b݉1p�`]�iA�y CV�zP �z�}x�}yu�8��	q�ypse����r57� Inp���xy͉576��(p+�)� ����|z� "Al�~w6\aYb����j8<�B؝�h ��PR<�J8��zPxC;�8�J�p�s��P��}x96\ {�(P|y�����A}x9 �� -��iv{�R� DM<�H7�zH-6�{66�3�1}x�[�tor�����P��y�m�!��sZ��]�2����naldۺ��)�޸stK���}str��ypsk��=�\p����}x/j932|�C�� }�)}x8R}x2}���2��.|�޸_w���}hk_k�FH��z9!�}xke*�n�95�
���yhe�z@sk�,�f�l.��H�et_w|y�"}yac� �y� �zbak��H�Z�ent��h�\	m���s���� � �d�༛�Y�;�(�Z�(�@�z9Pf|yv�@�� .������ l�n�( Ll�gd��=
i���! Z���+�00iB\�H[�H���� z-�h[�C" #���82��2�@}�ORp��� ���iB/̿LN@�"F���f���h@+�=���t{z OR����83�i1�3t ˚�~nc+���fc����5���8�35�z����i�;�5�:�B�ri��ER����b݉ (ˊngQ,�@�,4�*R0ȭY�k��mo�`]/r��p�+��ptp�z(�5\pk�=O?��� �0[ڈ��0�/�/ ?S�i�k߽�ij��
���?�+�db��� s50l�a��x���S�[d G�yϋ�cce��0K�50�Kz1|y�6��J�e�RDE��y|A;nt�
 Pa��(��9\g{�H�919�[�END�\:� V=i��tool<?ވ:	�J[�uppK/=_��vk{��K[��Z� �Z��O�O�O�8�OK�8H��?�_rj;*h��ndr{�H]end$��Ir:�(�3��o�~H73;���/�&7 ;*��{X�j�|����"�4�  am_x�O�ve�ʘ���v$I���o�?|�xj{���� �Tz{�] R�5;�J9�;989@ﭹ���_��p�m
��
�`����e�kR� R�}++R7�J L:;) "���KzR�/p+zx�d	�-��|�	�633�06� S�I~R6�sqt�z��:�LND��7IF K�45��-con{
C9�i�*�ar �jyp�	�d�s "����EN�l�y��s��l�gr括e-����8568��`�zrpi{�x=�H�4 l�^�wnj�! r˛vv�:�nn�}RC:| ��� J9�Z����8[67�13J;6���8 �JT�`(iR��R|"ٟc  STD���.pLANG(&�����r��ti�����P��q��)0-�� =E��kg
��y`� ��5����R73�0��(��8 (i^��ErrP��,�`���PC��x���rv�ge������8���g�e��a<����	�.ޠ�isio��ck#in�� �R�(���pGi� ������؁��j	��PFK�"��XA��\@��B�P4��!��d��agabbPbbb������P��P��(1��S�P�Р�FS J���J91��685b9!	��02*-4<627���Y��,����X�v��s\�GFSO8����sex��/�vr�����&��v�RG(R68'64����#8	�G (� CCR���I���cc�� �"CkH���9�\�RBT}rgOPTN�4�4�2��4�?�?O"Ocrg�.8EF��DP)N����
hEd�iD�ion hEnd.qhExa�FINThER��7hE� nhEa�@�hE�0"hEHQhEhd\m�FHD�F�iD\erh�F���O�A�ihE��sF�"Uir�ehEhiDtiDrh �@�tdB�t��t��tn An�_��j0�tt2�t8�t0E�t�a�U�`t f�1�t�2�t� m�U�a�U葈U-`As�U�ѠW
 �t1�ލt�6��U R�88�U851_f4<�`�Utiar�U���tit� �tl"�tM�R S�f`�fTX�P�U��epm�f"w #1�f! T�fy��fm�g��e�P�U� 2�U 70�Uon�jg�t�@_f J7r�Vipp�fon,�U����X�v4m�j79b�fc��e]h98jg��"m�\chp�WE�N�vd@Pb{StoD'�� E f�@�VgF0��el�gxшU��jA8svY��f�m�6uh�arel�UKARNo�Comc�u�RĆeL*wp\ �V
+v�Y�u�fp\e�VA�N"���k�gpcp_f1a!I�[�f4y��wf
! Gf C�o�uarwf�FvІ84_f5 H�f�H84�v63 Hv�fH7�v779_fi24��7rw69*�+65�f1�g8p��V�75�VIC �f ;AP7v893���0R0m��B�eck���Hs�
E����#fMNS+v�ПVՐ�V�P_f-]�_�Q�VX�\���tch믅ԈUw3\pSfWT"_f��_�_hin_� �0�3jgoX�е(ROB�wOG���AUe�A �^�HR�PxflR�uuyQuug_Sf̉3nuh523�Vle*wOrity �6�2��6�5sv54f�4�І40����H60b�v0�h�[�08�@�+�=�O�a���8< ���68v�`��s�C75^0��A�rw7�Рh����וл�3�v3�Y� е ��େ2f���� 2�9#f�p���\ib<f��;sbs�w��oG scbP1oCja��Ly2%� -k�E"��74�9 wf (W�_�	`��XPF���w�vF�E�X�Ϯ`wep�Vp��a\wvTf�͸�z50+�"WV����֤u��2�Y �� ��nte�g����^�f04 (�gx��8D����BPXk���!I/��`o�d�@���G��pv kϥ�ib�hp
om ��wfE�A�f��Hfdn���z8Z�f�_�F�Vra�W�_�oi �v<�al�VVAx�V��2�� 996#fV�CA��,�vast�#/�q� ��"�dp6/fyn:�fi����58����D��odcif��.e8DP��tq (d��o "�� �o��Rg�d9Ԑ'G���strS���OAW����wR73�v16�"� Rf�79�2\���iTra��c�ht�/�wv"TP+v\̀��tpe�c�w�or���+RC�59��8�� S5+�809�?��C�f�"�z\mߦD6�v��RE��$FL&�0�pcz�6�ve�rv�gng_��7�46�_��S_� Cqh�?�� �`%/@s�th��0�W897i3�g����m��f!��a$��x���� T������� ���rk�����`s�H�VAG�ǧset99����7��$F�EAT_ADD �?	����q�p��	x�� ����*�<�N�`� r���������̏ޏ�� ��&�8�J�\�n��� ������ȟڟ���� "�4�F�X�j�|����� ��į֯�����0� B�T�f�x��������� ҿ�����,�>�P� b�tφϘϪϼ����� ����(�:�L�^�p� �ߔߦ߸������� � �$�6�H�Z�l�~�� ������������ � 2�D�V�h�z������� ��������
.@ Rdv����� ��*<N` r������� //&/8/J/\/n/�/ �/�/�/�/�/�/�/? "?4?F?X?j?|?�?�?��tDEMO ^~�y   x �=�?�?OO%OROIO [O�OO�O�O�O�O�O �O__!_N_E_W_�_ {_�_�_�_�_�_�_o ooJoAoSo�owo�o �o�o�o�o�o F=O|s��� ������B�9� K�x�o�������ҏɏ ۏ����>�5�G�t� k�}�����Οşן� ���:�1�C�p�g�y� ����ʯ��ӯ ���	� 6�-�?�l�c�u����� ƿ��Ͽ����2�)� ;�h�_�qϋϕ��Ϲ� �������.�%�7�d� [�m߇ߑ߾ߵ����� ����*�!�3�`�W�i� ������������� &��/�\�S�e���� ������������" +XOa{��� ����'T K]w����� ��//#/P/G/Y/ s/}/�/�/�/�/�/�/ ???L?C?U?o?y? �?�?�?�?�?�?O	O OHO?OQOkOuO�O�O �O�O�O�O___D_ ;_M_g_q_�_�_�_�_ �_�_
ooo@o7oIo como�o�o�o�o�o�o �o<3E_i �������� �8�/�A�[�e����� ��ȏ��я�����4� +�=�W�a�������ğ ��͟����0�'�9� S�]�����������ɯ �����,�#�5�O�Y� ��}�������ſ�� ��(��1�K�Uς�y� �ϸϯ���������$� �-�G�Q�~�u߇ߴ� �߽������� ��)� C�M�z�q����� ��������%�?�I� v�m������������ ��!;Eri {������ 7Anew� �����/// 3/=/j/a/s/�/�/�/ �/�/�/???/?9? f?]?o?�?�?�?�?�? �?O�?O+O5ObOYO kO�O�O�O�O�O�O_ �O_'_1_^_U_g_�_ �_�_�_�_�_ o�_	o #o-oZoQoco�o�o�o �o�o�o�o�o) VM_����� �����%�R�I� [����������Ǐ� ����!�N�E�W��� {�������ß���� ��J�A�S���w��� ������������ F�=�O�|�s������� ���߿���B�9� K�x�oρϮϥϷ��� ������>�5�G�t� k�}ߪߡ߳������� ��:�1�C�p�g�y� ������������	� 6�-�?�l�c�u����� ����������2) ;h_q���� ���.%7d [m������ ��*/!/3/`/W/i/ �/�/�/�/�/�/�/�/ &??/?\?S?e?�?�? �?�?�?�?�?�?"OO +OXOOOaO�O�O�O�O �O�O�O�O__'_T_ K_]_�_�_�_�_�_�_ �_�_oo#oPoGoYo �o}o�o�o�o�o�o�o LCU�y �������	� �H�?�Q�~�u����� ����׏����D� ;�M�z�q��������� ӟݟ
���@�7�I� v�m��������ϯٯ ����<�3�E�r�i��{�����˽  ¸����)�;� M�_�qσϕϧϹ��� ������%�7�I�[� m�ߑߣߵ������� ���!�3�E�W�i�{� ������������� �/�A�S�e�w����� ����������+ =Oas���� ���'9K ]o������ ��/#/5/G/Y/k/ }/�/�/�/�/�/�/�/ ??1?C?U?g?y?�? �?�?�?�?�?�?	OO -O?OQOcOuO�O�O�O �O�O�O�O__)_;_ M___q_�_�_�_�_�_ �_�_oo%o7oIo[o moo�o�o�o�o�o�o �o!3EWi{ �������� �/�A�S�e�w����� ����я�����+� =�O�a�s��������� ͟ߟ���'�9�K� ]�o���������ɯۯ ����#�5�G�Y�k� }�������ſ׿��� ��1�C�U�g�yϋ� �ϯ���������	�� -�?�Q�c�u߇ߙ߫� ����������)�;� M�_�q������� ������%�7�I�[� m�������������� ��!3EWi{ ������� /ASew�� �����//+/ =/O/a/s/�/�/�/�/ �/�/�/??'?9?K?�]?o?�?�?�?�?�9  �8�1�?�? 	OO-O?OQOcOuO�O �O�O�O�O�O�O__ )_;_M___q_�_�_�_ �_�_�_�_oo%o7o Io[omoo�o�o�o�o �o�o�o!3EW i{������ ���/�A�S�e�w� ��������я���� �+�=�O�a�s����� ����͟ߟ���'� 9�K�]�o��������� ɯۯ����#�5�G� Y�k�}�������ſ׿ �����1�C�U�g� yϋϝϯ��������� 	��-�?�Q�c�u߇� �߽߫��������� )�;�M�_�q���� ����������%�7� I�[�m���������� ������!3EW i{������ �/ASew �������/ /+/=/O/a/s/�/�/ �/�/�/�/�/??'? 9?K?]?o?�?�?�?�? �?�?�?�?O#O5OGO YOkO}O�O�O�O�O�O �O�O__1_C_U_g_ y_�_�_�_�_�_�_�_ 	oo-o?oQocouo�o �o�o�o�o�o�o );M_q��� ������%�7� I�[�m��������Ǐ ُ����!�3�E�W� i�{�������ß՟� ����/�A�S�e�w� ��������ѯ���� �+�=�O�a�s����� ����Ϳ߿���'� 9�K�]�oρϓϥϷ� ���������#�5�G� Y�k�}ߏߡ߳����� ������1�C�U�g� y������������ 	��-�?�Q�c�u��� ������������ );M_q��� ����%7 I[m���� ���/!/3/E/W/ i/{/�/�/�/�/�/�/ �/??/?A?S?e?w?��?�?�?�?�1�0 �8�?�?OO1OCOUO gOyO�O�O�O�O�O�O �O	__-_?_Q_c_u_ �_�_�_�_�_�_�_o o)o;oMo_oqo�o�o �o�o�o�o�o% 7I[m��� �����!�3�E� W�i�{�������ÏՏ �����/�A�S�e� w���������џ��� ��+�=�O�a�s��� ������ͯ߯��� '�9�K�]�o������� ��ɿۿ����#�5� G�Y�k�}Ϗϡϳ��� ��������1�C�U� g�yߋߝ߯������� ��	��-�?�Q�c�u� ������������ �)�;�M�_�q����� ����������% 7I[m��� ����!3E Wi{����� ��////A/S/e/ w/�/�/�/�/�/�/�/ ??+?=?O?a?s?�? �?�?�?�?�?�?OO 'O9OKO]OoO�O�O�O �O�O�O�O�O_#_5_ G_Y_k_}_�_�_�_�_ �_�_�_oo1oCoUo goyo�o�o�o�o�o�o �o	-?Qcu �������� �)�;�M�_�q����� ����ˏݏ���%� 7�I�[�m�������� ǟٟ����!�3�E� W�i�{�������ïկ �����/�A�S�e��w���������ѹ�$�FEAT_DEM�OIN  ִ����ΰ�INWDEX�����ILECOMP �_���7����-�SET�UP2 `7��A��  N �l�*�_AP2BC�K 1a7� G �)Ҹ�ϯ�%�� ��&�:�����Ե��*� ��N���[߄�ߨ�7� ����m���&�8��� \��߀��!��E��� i������4���X�j� ��������S���w� ��B��f��s �+�O��� �>P�t�� 9�]���(/� L/�p/�//�/5/�/ �/k/ ?�/$?6?�/Z? �/~??�?�?C?�?g? �?O�?2O�?VOhO�? �OO�O�OQO�OuO
_ �O_@_�Od_�O�_�_ )_�_M_�_�_�_o�_ <oNo�_roo�o%o�o��oF�z�P~� 2>��*.VR�o�`* F�cLp�ZepPCx��`OFR6:��~\��{T��'��u��Q����w�Yf*.F
���a	�s��Ռ�d�����STM @�"�-��p�Y��`�iPendant PanelY���HO���?���[�����GIF�6�A��"�ߟ񟆯��JPG ����A���c�u�
��z#JS�=��`У+���%
JavaS�cripti���C�SZ���@���k� %�Cascadi�ng Style Sheets��_`
ARGNAMOE.DT�lD��\0��P�`�q��>`�DISP*g�JπD����σ����ϡ�	?PANEL1��O�%D�8�x�k�}�+�2m���b���~ߐ�%�0�3��W�b�E�����0�4u���b�������-�(�TPEIN�S.XML4���:�\H���Cust�om Toolb�ar����PASS�WORD��}nF�RS:\���� %�Passwor�d Config XoV��O��o� ?��u
�.@ �d��)�M �q�/�</�`/ r//�/%/�/�/[/�/ /?�/�/J?�/n?�/ g?�?3?�?W?�?�?�? "O�?FOXO�?|OO�O /OAO�OeO�O�O�O0_ �OT_�Ox_�__�_=_ �_�_s_o�_,o�_�_ bo�_�ooo�oKo�o oo�o:�o^p �o�#�GY�} ���H��l���� ��1�ƏU������ � ��D�ӏ�z�	���-� ��ԟc������.��� R��v������;�Я _�q����*���#�`� ﯄������I�޿m� �ϣ�8�ǿ\���� ��!϶�Eϯ���{�� ��4�F���j��ώߠ� /���S���w߉��� B���;�x���+��� ��a�����,���P� ��t�����9���]� ����(��L^������� �$F�ILE_DGBCK 1a��� ��� �( �)
SUMMARY.DG��hMD:�0�t Diag S?ummary1>
�
CONSLOG�&	t�CC�onsole l�og�=	TPA'CCN�/%�4/�?TP Acc?ountin�>
�FR6:IPKDMP.ZIPh/�l
�/�/@P Exception�/�n+MEMCHECCK*/�@?��Memory D�ataA?�LN?�)	FTP��?�'?�?K7�mme?nt TBD�?u7� >)ETHERNET�?f�!�OHOCEthe�rnet �fi�gura�/D�1DCSVRF�?�?�?��OQ1%�@ v�erify alyl�O�M,��EDIFF�O�O�OO_�R0%�Hdif�fQ_W�!�@CHG�D1F_-_?_�_ �f_�_S+P�Y2p�_�_�_Xo �_ooGD3No5oGo��o no�f�UPDATES.�"piFRS:�\ a}DUpd�ates Lis�tafPSRBW�LD.CM�h�Lr�c�PS_R?OBOWEL�?<}�aHADOW�o�o�of�Q3Sha�dow Chan�gesi��==�&�NOTI�OA��S��O5Noti�ficqB���O�AJ?�nc��p� ��D��L��󟂟� ��;�M�ܟq� ����� 6�˯Z��~���%��� I�دm�����2�ǿ ٿh�����!�3�¿W� �{�
ψϱ�@���d� ��ߚ�/߾�S�e��� ��߭߿�N���r�� ���=���a��߅�� &��J��������� 9�K���o����"��� ��X���|�#��G ��k}�0�� f���,U� y��>�b� 	/�-/�Q/c/��/ /�/:/�/�/p/?�/ )?;?�/_?�/�?�?$? �?H?�?�?~?O�?7O �?DOmO�?�O O�O�O VO�OzO_!_�OE_�O�i_{_�$FILE�_LpPR[p���_P�����XMDONLY� 1a�UZP 
 �
_�_._oR_ o;o__o�_�o�o$o �oHo�o�o~o�o7 I�om�o� �� V�z�!��E�� i�{�
���.�ÏՏd� �������*�S��w� �����<�џ`���� ��+���O�a�🅯�੯8���߯�ZVIS�BCK�X�Q�S*�.VD�0���F�R:\��ION\�DATA\�â���Vision� VD file \�j�����̯ڿį�� ���4�ÿX��|ώ� ϲ�A���e�w�ߛ� 0�B���f��ϊ�ߛ� ��O���s����>� ��b�����'���� ��������'�L��� p������5���Y����}���$�ZMR2_�GRP 1b�[��C4  B� 	 �Qk}h �E�� E�  �F@ F�5U��/
h L���M���Jk�K��v�H�,�H�k��?�  x�/h 9tQv�8���6h�%<�A�  3E�BHeB�a `�E@i/g��^h @UUU�U���>�]�>П��;r8	=�==E��<D��><�ɳ<��Ε�:�b�:�/'79�W�9�
@�8�8�9��T/�Q/�/�eE7� E?p� D�D�/�D��  D�  C���/9
_CFG =c�[T �/?�0?B?�NO ^�Z
F0x1 }0��RM_CHKT_YP  �P� h�P�P�P��1OM�0�_MIN�0
����0�PX�PSSuB�#d�U�Pi�?	�3O$O�U�TP_DEF_O�W�P
�Y?AIR�COM�0JO�$G�ENOVRD_D�O�6�RxLTHRֺ6 d�Ed}D_E�NBiO }@RA�VCGe�7� ���FnH E��� Ga H��� H�@JCh`�/O?_�G_�X_{ ��AOUZ�@kN {<NB{8���_�y_�_�_�_  C�
a �a �%o�?doCOm?aUc~	�Y+O.�@SMT�Cl�IZ ��04d�$HOST�C�"1m�Э 	
x
{�
:bye V�����zu�� ��$�GH��p	a�nonymous K�y���������	 -�A�c�V�h� z������ԟ��� �M�_�@�R�d�v��� ˏݏ����7�� *�<�N�`��������� ��̿�!�3��&�8� J�\ϟ���ïկ׿�� ������"�4�w�X� j�|ߎߠ�������� ����0�sυϗϩ� �ߜ������������ K�,�>�P�b���s��� ����������G�Y� k�L�p���� ��� $6Y Z��~����	 �-? /SuB/h/ z/�/�/��/�/�/�/ 
?-/_qR?d?v?�? �?��//?�?I/ *O<ONO`OrO�/�O�O �O�O�OO3?E?&_8_�J_\_n_�g�aENT� 1n�i�  sP!�O�_  �@�_�_�_o�_+o�_ Ooo[o6o�o�olo�o �o�o�o�o9�o o2�V�z�� ���5��Y��}� @�v�����׏������ ��+��T�y�<��� `�����埨�	�̟ޟ�?��c�&���J�QUICC0��p���㯦�1���ү3����24��"���!ROUTER��`�r��ӿ!PCJOG�Կ��!192�.168.0.1�0����CAMPRYT$� �!�1�K�2�RT��O�a�����TNAME !~�Z!ROBO=����S_CFG 1�m�Y ��Auto-st�arted�4FTP�?[��?�O�� O�߼������ߋO� (�:�L�o�]����0�������#��:4� F�X�9�l��P����� ����z�������# F���Yk}��� �?�?�?�?.b�C Ugy�N��� ���-/?/Q/c/ u/�/��� /�/ 6?)?;?M?_?"/�? �?�?�?�?�/p?OO %O7OIO[O�/�/�/tO �?�O
?�O�O_!_3_ �?W_i_{_�_�O�_D_ �_�_�_oo/orO�O �Owo�_�o�O�o�o�o �o�_+=Oa�o ������4o FoXojoK�~�o���� ����ɏ�����#� 5�X�ڏk�}������� ş��,�>�@�1�t� U�g�y�����`���ӯ ���	�,���?�Q�c��u�������_ERR� o�ʡ���PDUSIZ  3��^L��ȴ>�W�RD ?"����  guest-�!�3�E�W��i�{���SCDMN�GRP 2p"�;˰��3���-�K�� 	P01.05 8��� �����>,�j�  2�1�� ~� ���T����������_�����$���`ϿQ�<�u�`�������  �o  
��N(��P,�(����Qo���������kl�� 8�#{��d�����"ߙ�_GWROU��q�������	����4S�Q?UPD  �ȵYX��TY������TTP_AU�TH 1r�� �<!iPend�an����8�g��!KAREL:q*����KC-��=�O�%�VISI?ON SETb����3�#�������"�  ��_6H��l~��CTRL �s�����3���FFF9E3���FRS:DE�FAULT�FANUC We�b Server ����	�Ĵ}�������WR_�CONFIG �t�� ��I�DL_CPU_P5C*3�B��I w BH/%MIN:,���M%GNR_IOັ���Ƿ1 NPT_SIM_DO&��+STAL_S�CRN& ��*T�PMODNTOL8�'�+bRTY�(I!8�&����ENB�'���-$OLNK 1u���Q?c?u?�?�?�?�?52MAST�E~ ��52SLAV�E v��34��O�_CFG�?IUO���OBCYCLE�>OD$_ASG s1w����
 �? �O�O�O�O�O�O__ 1_C_U_g_y_�_�;tBWNUM�Ĺ
B�IPCH[O��@R?TRY_CN*�"@ĺB�!���P1�ȵ1 B;@Bx�>��Jo�1 SDT_I�SOLC  ���f��$J23_D�S4�:��`OB�PROC?�%JOmG^�1y�;��d8�?��[D�o�_?؟֟O|QN s��V����-�~o�h�`Y A�_>�bPOSRE�o�&?KANJI_�0����/k�+�MON zg��2�y�Ϗ�@���Ҿ)�0c{,��9�T�f�CL_�LY �R�_k�EYL_OGGIN@�����ȵ�$LA�NGUAGE �k2ENGL�ISH 㑱�LG�1b|�2���3�x������O � {'0,�� �
q��3�MC:�\RSCH\00�\��LN_DI�SP }�?f��MKm�OC�"@"D�zh#�A�OGB?OOK ~K��`w���w�w���X�� �-�?�Q�c�u���11����	����h�޿����ॐ_B�UFF 1@=���)�����E� a�sϠϗϩ����� �����B�9�K�]߀oߜߓߥ��ߜ��D�CS �� =��͗�ֿM�l:��L�^�p���IO 1�K No�� ����������� %�9�I�[�m������� ����������!3hEY��Ex TMlnd������ 0BTfx�� �����//��N�SEV`}��TYPln��/�/�/)-P�RS�P���>bFL 1���`��?,?>?P?b?t?�?�/TP��loq"}��NGNAM�d���Ւ��UPSu�G�I�U\�e�1_L�OAD�`G %�}�%REQME�NU�?�\MAXUALRM�Wk�X\@N�1_PR�T`ԣ4��Z@Cx��ꩦ���OV�9ŜC�`P 2]��K �9�	q!�P]  � �OQ�R9_$_6_o_� ]_�_�_�_�_�_�_�_ oo@oRo5ovoao�o }o�o�o�o�o�o* N9rUg�� �����&��J� -�?���k�����ȏڏ �����"���X�C� |�g�������֟���� ݟ�0��T�?�x��� m�����ү��ǯ�� ,��P�b�E���q����SGD_LDXDI�SA�0�;��MEM�O_AP�0E ?=�;
 j �� ��*�<�N�`�rτ�~Z@ISC 1��; �����T�A����ϛ�$��Hߙ�C_MSTR �B-~g�SCD 1����<߶�8��������� "���X�C�|�g�� ������������	� B�-�f�Q���u����� ��������,< bM�q���� ���(L7p [������ /�6/!/Z/E/W/�/ {/�/�/�/�/�/�/? 2??V?A?z?e?�?�?��?X�MKCFG ��vݽO�CLTAWRM_�2��G�B� P�2�@>OFD{@M�ETPU�C�@���~�ND�@ADCO�L`E�@kNCMNT�O tEo� ��v��N5C.A�O�DtEP�OSCF�G�NPgRPM�OYST@{1��� 4@��<#�
oQ�1oU_ �Wk_�_�_�_�_�_�_ o�_oOo1oCo�ogo�yo�o�o�o�o�atAS�ING_CHK � �O$MODA�QC��?���>+uD�EV 	��	�MC:_|HSIZ�Eѽ���+uTAS�K %��%$1�23456789� ��u)wTRIGW 1���l#E%�̀)����S�6�%C�vY�P�q>�At*sEM_INF 1�#G� `)�AT&FV0E�0`�׍)��E0�V1&A3&B1�&D2&S0&C�1S0=ƍ)A#TZ׏+��H/�W��K���A����j�ӟ����	� ��.�� �����;����Я ⯕����*�<�#�`� �%���I�[�m�޿� ���K�8����n�)� ��y϶���{��ϟ��� ÿտF���jߡ�{ߠ� S������������� ��T���+ߜ��a� ��	�����,���P� 7�t���9��]�o�� ����(:q�^���=����XN�ITOR�@G ?�s{   	EOXEC1�32%3%4%5%�p'U7%8%9�3  ��$�0�<� H�T�`�l�Px���2�2�U2�2�2�2�U2�2�2�2��3�3�30+qR�_GRP_SV ;1��� (�?�/�'u�q_D{�~�1P�L_NAME �!#E0�!D�efault P�ersonali�ty (from� FD) �4RR�2�! 1�L6�8L@�1P
d d�/v?�?�?�? �?�?�?�?OO*O<O NO`OrO�O�O�O�O�O�OJx2e?_ _2_D_�V_h_z_�_�_�_r< �O�_�_�_o"o4oFo�Xojo|o�o�o�i�VD�_�n
�o�oNtP�o *<N`r��� ������&�8� n���������ȏ ڏ����"�4�F�X� j�|�K�]���ğ֟� ����0�B�T�f�x����������Ү �FnH F�� gG=��'�"�����"d�$/�A�&� d�r��׭Ҫ�/����ٿܧ ͸���  ��0�6�T�v�̰��ϩ̾`A�   ��˿��Ǹ]0���ƿ 3�¿W�B�{ߍ�x߱�dB5K3�9^0`�!0 � ��0�� @D�  &��?����?� ��!A�����$���(;�	l�	 ���p�V� ]0M� � _� � �l�r����K(��K(��K ��J�n��J�^J&Ǔ�2���������@Y�,@Cz?@I�@���������N�����f���_�I_���SѬ�Ä���  <��% ß3������!?s8y�
�/�!��x����T� ܌�������}���    �������  ���������	'� � 0�I� �  ������:�È~TÈ=���l 	�(|�����ш����ψ��N<@0�  '����@2��@����@!����@)���C@0C��\C�I�CM�CQ�� ���ģ�%%����� ��B���@0��lc@� ��!Dz�߀�V�//+/Q/<"?�� �H@q)lq�%  �����  � p�!?��ff���/�/V/ ���/;=!8� !?/:@��D4�� \6Pf8`�)c�\�\��?Lv ��$<!;�Cd;��pf<߈<���.<p��<�?L:��ݧA����d����?fff�?�?&@��@��� B�N�@T�,E�	��	A�� �dO�O�7H��/�O �O�O�O _�O$__H_`Z_E_~_�MEF� m_�_i_�_UO�_yI�_t2o�XC��E��"?Gd G;ML!o �omo�o�o�o�o�o�o �o$H��iww9 ��_�o�U��*�<�ڪ����/�6�������ď��菎�AB�A�����C؏0=�ԏ��X��񨑟�,�����  �P��"@�<��E� AC���s��x�؄��(�����/�B�/�B"�}A��#�A��9@�dZ�?vȴ,��~�����<)�+�� =�G��j����q���
AC�
=C������년� ��p��Cc�¥��B=���f�f�{,�I����HD-�H��d@I�^�F8�$ D;ޓܪ����Jj��I���G�FP<����QpJnP�H�?�I�q�?F.� D��Ɵ g�R���v�������� п	���-��Q�<�N� ��rϫϖ��Ϻ����� �)��M�8�q�\ߕ� �߹ߤ߶�������� 7�"�[�F�k��|�� ����������!��� W�B�{�f��������� ������A,e P�t����� �+;aL��p�����(���g�3:��1��%�3�V��/"��(/:/�!4M㇬T/f/F1�=�Ӏ/�/4Ue'��T9�-�)�/�/?P�/4?"<]�P�2Pf>�q��?��?�?�?<�?�9���(�?�?�/OO?OeOPO�QB� hOzO�O�O�O�O�O�?`t.__R_@[/X_�b_�_�_�_�_�_�Q{f�_�_o
o@o.odo�rj  2 Fn�H"�F��"�G=b��B# ��C9)��@|�@��o�o�o �E�� F��`�H C����6E{�c��kE��q�da �O����{?ސ�q* ��D  zqu `�
 � !�3�E�W�i�{����� ��ÏՏ�������q� ��P+�~Y���$MSKCFM�AP  �%� ^f�q�q�p�D�ONREL  X5[��0D�EXCFENB��q
Y����FNC�����JOGOVLI�M��d����dD�K�EY�����_�PAN����D�R�UN��SFSPDTYw0�������SIGN����T1�MOT럜�D�_�CE_GRP 1-��%[�\�O� �O�&��d�Q��u� ,�j���b�Ͽ��Ŀ� ��)�;��_�σϕ� LϹ�pϲ��Ϧ��%� �I� �m��fߣ�Ov�D�QZ_EDIT���U��TCOM_�CFG 1�Q������"�
��_A�RC_��X5ؙT�_MN_MODE���縙UAP_�CPLF４NOCHECK ?Q� W5�H���� ������'�9�K�]��o�����������v�N�O_WAIT_L؉��׾�NT����Q��{_ERR�ȡ2�Q��1�  ��t���H*������`�OI�Px�  8%��!8�?nw�s5V�
BPARAM:J�Q���v	���7so� =�`3�45678901 �/ *�?/Q/-/]/��/�/u/�/�/�+�7��?<�7?��UM_RSPACEN��'2$�p?z4�$OD�RDSPE㌦��O�FFSET_CAqR�Ќ�6DIS�?��2PEN_FIL�E�0�$��֌1PT?ION_IO
���@M_PRG %\:%$*IO[N�3WORK �Χ=�� ���F7�"�Bh���@(7�A�	 ��x�C7��c���0RG_DSBOL  \5���|�_�1RIENTT5O��9�C��pZ���a�0UT_SIM�_DGX�+��0V~�0LCT �%��ҟDx=gT_PEX�h��?�TRATh� �d���T�0UP S�u^�Ӡ�o�o�_:oHi�$�2�ǣ�L68L�@�_S
d d '?�o�o�o�o�o�o�o 1CUgy��������I2 ~o'�9�K�]�o���������ɏ9�<��� �)�;�M�_�q����� ����H�j3�H1`��XRP�C�U�g� y���������ӯ��� 	��-�?�Q� �2��� ������Ͽ���� )�;�M�_�qσϕ�d� v���������%�7� I�[�m�ߑߣߵ���0��X���'��*��S%4H�Z�?�}������&?������ �@�����+�I�O��m�����?@������A�  ������� ���M8q\�@���z�d`O�P�1�k�ۆ�sd`�R0 ��D$@ @D��  DD?QD	��U��  ;�	l1	� ��p��s��j Կ � � ʉ���� H<zH<�W�H3k7G��CG���G9|+c	�H
���� +CC9P/9P49S;Q�9/��9  ·�  1!�H7 3����/1/C/��BY����>XQ�^�H�<Pq/ ܩ/�"2�#�3��.�   � �0�� �  0�6�/?��%	'� � �M2I� � � ���
=��a�q?�;�#&�(�3@�/�'�A�?4;�B�?�'NEPO  '�VP3D�b CEPC�W�\Cf Cj Cn/�@OROߑ  �����D%%~��� ��'�B���FEP�E˜@XP�E5z�_s/8_�#_H_n_�"�� ��H]2�Y�A�U M �C�H�A�0=p�Q?�ff���_�_s_ ��o(kZQ8�0>oLj-�!ad�'�0yfP�h�Y�yy��3?L�0�T�!;��Cd;�pf<�߈<��.<p��<�?ij��WA�Eل1d�31���?fff?�@?&�+p�$@��=r�?N�@T�IuՉ ��&q-ZP!�� we o����� �A�,�e�w�b����� ��я����l���tO��CE���2?Gd G;�|>� ����ß���ҟ��� �A�,�e�����V� ���د6���r�#�5�G�Y��Z� �_�f��������̿Ϡ&AB @A�@%���5�C���Z���/i�?����Ϗ��ϳ�U�P���2]!YNE� !CU%�̣�Ŀ�����E�@I�!t�B��/B"�}A���#A��9@��dZ?vȖ+����~��<)�+� =�G�(���Ԁ�q���
�AC
=C������녡� ���p�Cc�����B=���ff�{���I���HD-��H�d@I�^�?F8$ D;������̠Jj��I��G�F�P<��QpJn�PH�?�I��q�F.� D� �E�τ�o������ �����&��J�5�n� Y�k������������� �� F1jU� y������ 0T?xc�� �����//>/ )/;/t/_/�/�/�/�/ �/�/�/??:?%?^? I?�?m?�?�?�?�?�?  O�?$OOHO3OXO~O�iO�O�O�O�O�O��(�}���3:�O�a�y�)U�E3�V�_+_9R�E_W_t��4M��q_�_t���=ӝ_�_4Ue'��T9�]�Y	o@�_-ooQo?lz�P�b	P�n�����o�O�o��o�o�i���( L7\�mt�B����������o��K�9�o�]�/u������ŏ�ُ�{f��9�'�]��K�����  2 wFnH��F�Щ֋G=��B@P!�.�C9F��p��@2���	���C�E�� F�>���H C���S�b�����������¯ԯ��?����Jy�C�C�|�C�}�
 ۯ>�P� b�t���������ο�����(ϧ�� ���m[�~Y��$�PARAM_ME�NU ?�U��  �DEFPULS�E4�	WAIT�TMOUT��R�CV�� SH�ELL_WRK.�$CUR_STY�L����OPT����PTB����C���R_DECSN ��teG�A�S�eߎ߉� �߭������������+�=�f�a�SSREL_ID  �U��a�u�USE_P�ROG %p�%8b���v�CCR������ax���_HOST7 !p�!������T�`��8�����:�t���_TIME����a�GDE�BUG��p�v�GI�NP_FLMSK̝���TR����PG�A�� ��{�CyH����TYPEm�y�a�[��� ���!JE Wi������ ��"////A/j/e/ w/�/�/�/�/�/�/�/�??B?��WORD� ?	p�
 	�RS��sPNeSu��~2JO��rTE[��?CCOLu>8�?>L�� �P��p���T�RACECTL �1��Uz� ��`��)O3BFD/T Q��U^@#@�D � sckO}O�O�O�O�O�O �O�O__1_C_U_g_ y_�_�_�_�_�_�_�_ 	oo-o?oQocouo�o �o�o�o�o�o�o );M_q��� ������%�7� I�[�m��������Ǐ ُ����!�3�E�W� i�{�������ß՟� ����/�A�S�e�w� ����gO��ǯٯ��� �!�3�E�W�i�{��� ����ÿտ����� /�A�S�e�wωϛϭ� ����������+�=� O�a�s߅ߗߩ߻��� ������'�9�K�]� o����������� ���#�5�G�Y�k�}� �������������� 1CUgy�� ������	- ?Qcu���� ���//)/;/M/ _/q/�/�/�/�/�/�/ �/??%?7?I?[?m? ?�?�?�?�?�?�?�? O!O3OEOWOiO{O�O �O�O�O�O�O�O__ /_A_S_e_w_�_�_�_ �_�_�_�_oo+o=o Ooaoso�o�o�o�o�o �o�o�9K] o������� ��#�5�G�Y�k�}� ������ŏ׏���� �1�C�U�g�y����� ����ӟ���	��-� ?�Q�c�u��������� ϯ����)�;�M� _�q���������˿ݿ ���%�7�I�[�m� ϑϣϵ�����������!�3�E�W�a��$�PGTRACEL�EN  b�  ��a���w�_UP �/������В��  ��w�_CFG7 �����a�����������������DEFSP/D ���`щ���w�IN��TROL �����8��F�PE_CONF�I�Ш���������LID�ө��	��LLB� 1��� �t�B� � B4��� ���� ���� 8?8�?�0�K� 0�G�i�k�}������� ������5Ak�����2���	�?��GRoP 1���lb��A�  �333�a�A��D�@� D�� D@� A@�Ta�d�+������� a	='����´#��B 9!///�O/9/s/
��?�����/�/�.�/ �=o=	7L �/?�/?P?;?t?_?��/�?�??�?�?�? G DzC Oa�
O HO�?XO~OiO�O�O�O �O�O�O_�O_D_/_�h_S_�_�Z!a�
�V7.10bet�a1�� Ax;���R��y�Q�?���Q>�\�)�QB0���PA���SBp���QA�9Sy�b
a�S ��_2oDoVoho��Ap���"���o�o�o�o��ة�KNOW_M�  ��֦�SV� ������5O8J\u_�@k}��Ҵ��M]��z�Д�R	��%%�"��|~���� ��u��P@�a�]�a�q�Xm��Ц�MR]��} ��&%O�P�$ӏ�K{ST]1 1���
 4��vi�Q:� �"�4�F�w�j�|��� ����ğ	����?�� 0�u�T�f��������P��ү��2� ��a��<K��^3 5�G�Y�k��4���������5ۿ���ς�6.�@�R�d��7 �ϓϥϷ��8�������
��MAD  ����)�OVL/D  ��G��PARNUM � ������T_S+CHy� ��
���8��0�UPD���������_CMP_0�p|�pp'�e��ER_CHK������j����RS8��oW_MO{����_���_RES_G��� o��� ������������ 2%VIzm`�R�4�\�l��Q���� ��S�ڰ�S� -�9X]S��x� �S������S�&���//S�V 1����a�q@c?\��THR_INRЮ�~��r�ed�&MA�SS�/ Z�'MN��/�#MON_QU?EUE ���fT"��a��N��U��qN�&��0END1;�79EXEF?75\��BEE0'?3OPT�IO$7D�0PROGRAM %�*�%0T/��2TA�SK_I{ԍ>OCFG ��/���?^"@DATA�s�+K��"�2��O�O �O�O�O�O�O_!_3_�E_�Oi_{_�_�_ROIWNFO�s�oM�
4 [_�_
oo.o@oRodo vo�o�o�o�o�o�o�o *<N`�W�T��oL �	!A�K�_%A�+I�^�vECNB|б}���v2���xG%A2��{ �P(O�4�F� �C�e��z_EDIT �+O����>DWERFLg8|#� �RGADJ M��:A����?"���!߆1�q�]�?�?���A<@��v%<�l�ӈ����q2�)��R	�H0le�{"6�?�
��AF$�t$�ܖ*�/� **:��"����� d�1�f�Ցd�[�B U�#���3�E�s�i�{� ������߯կ�a�� �K�A�S�Ϳw����� ����9����#��+� ��O�aϏυϗ�߻� �������}�'�9�g� ]�o��ߓߥ������� U����?�5�G���k� }����-������ ����C�U���y��� ����������q -[Qc���� ��I�3);��_q���t&	 >O@/Հ./g/R$ݙ�/�ߓU/�/Q/�/�/�P?REF �)�Հ�Հ
߅IORI�TY�72F��MP�DSP�1яG7UT�FǓކODUCT�
A�:�/��OG��_TG΀B����2TOENT 1�� (!AF_INEq0OG?!tcpO6M�!ud%O^N!icmMOu��2kXY"�Í��X1�)� ��O�OX0��O�O�E�O)__M_ 4_F_�_j_�_�_�_�_ �_o�_%o7o*�3"���=Y�yo�o��>�+�J��/�io��o�������AK�,  �0�q'�9K]X5�7�pHA?NCE �)��rrn{d�o��uyw	3��?"3ق�POR_T_NUMr3X0����_CAR�TREPR0����SoKSTAq7 C��LGS @ȍ���K�X0Unothing�����̏�܌�����#��?k�T?EMP ɕ94�����_a_seiban�/���/�� ͟���ܟ� �9�$� ]�H�Z���~�����ۯ Ư����5� �Y�D� }�h�����ſ��¿�� ��
�C�.�g�R�w� �ψ��Ϭ�����	��� -��*�c�N߇�r߫� ���ߺ������)��M�8�q�\��6�k�VOERSIP0�7��� disab�le�r<�SAVE� ʕ:	26�00H844����,�!�.�@�_Od�C 	��{2 /����X�e����	-;
��c�n ��L��]_�0 1˧K�� "����0/URGE�pB�0T6l>5�WF� DOr6��r�6W�0�"�W�RUP_DELA�Y �;�R_?HOT %%&~1���+R_NORMALy�2���SEMI��"/�!_QSKIP���w�x��g/��/�/�/ r-�5�/�'�/??(? �/L?:?\?�?�?�?l? �?�?�? OO�?"OHO 6OlO~O�OVO�O�O�O �O�O_�O2_ _V_h_ z_@_�_�_�_�_�_�_����$RBTIF�?�RCVTMO�UT�B��`D�CR��E) ��~!-�1�C����C���A�7�f�/|/ ��?�$�a9�o�o��o ;�Cd;��pf<߈<���.>�]�>П��o��o'8} 8^p�� ����� ��$��1%RDIO_TYPE  �.��EFPOS1 1}���  x�� ���Ώ���{�� ��:�Տ7�p����/� ��S�ܟ���՟6� !�Z���~����=��� دs����� ���D�V� ��=�����¿]�� ��
ϥ��@�ۿd��� ��#ϬϾ�Y�kϥ�� ��*���N���r��o� ��C���g��ߋ��&� �����n�Y��-�� Q���u������4��� X���|���)�;�u��� ��������B��? x�7�[�� ���>)b�� !�E��{/� (/�L/^/�/E/�/ �/�/e/�/�/?�/? H?�/l??�?+?�?�? a?s?�?O�?2O�?VO �?zOOwO�OKO�OoO �O�O_._�O�O_v_ a_�_5_�_Y_�_}_�_ o�_<o�_`o�_�o�o|�2 1ш�2oDo ~o�o�o &oD�oh e�9�]�� 
�����d�O��� #���G�Џk�͏��� *�ŏN��r���1� k�̟��🋟���8� ӟ5�n�	���-���Q� گu�����ӯ4��X� �|����;���ֿq� ����Ϲ�B�ݿ�� ;Ϝχ���[����� ���>���b��φ�!� ��E�W�iߣ����(� ��L���p��m��A� ��e���������� �l�W���+���O��� s�����2��V�� z'9s��� ��@�=v �5�Y�}�� �</'/`/��//�/ C/�/�/y/?�/&?�/ J?�/�/	?C?�?�?�? c?�?�?O�?OFO�?�jOO�O)O�O�o�d3 1ҵo_OqO�O)_ _M_SOq__�_0_�_ �_f_�_�_o�_7o�_ �_�_0o�o|o�oPo�o to�o�o�o3�oW�o {�:L^�� ���A��e� �b� ��6���Z��~���� ��Ə �a�L��� ��� D�͟h�ʟ���'� K��o�
��.�h�ɯ �������5�Я2� k����*���N�׿r� ����п1��U��y� ϝ�8Ϛ���n��ϒ� ߶�?�������8ߙ� �߽�X���|���� ;���_��߃���B� T�f�����%���I� ��m��j���>���b� ����������i T�(�L�p� �/�S�w $6p����/ �=/�:/s//�/2/�/V/�/�O�D4 1��O�/�/�/V?A?z? �/�?9?�?]?�?�?�? O�?@O�?dO�?O#O ]O�O�O�O}O_�O*_ �O'_`_�O�__�_C_ �_g_y_�_�_&ooJo �_no	o�o-o�o�oco �o�o�o4�o�o�o -�y�M�q� ��0��T��x�� ��7�I�[������� ��>�ُb���_���3� ��W���{������ß ��^�I������A�ʯ e�ǯ ���$���H�� l���+�e�ƿ��� ��ϩ�2�Ϳ/�h�� ��'ϰ�K���oρϓ� ��.��R���v�ߚ� 5ߗ���k��ߏ��� <�������5���� U���y������8��� \�������?�Q�c� ������"��F��j g�;�_��x�/45 1�? ���n��� f���%/�I/� m//�/,/>/P/�/�/ �/?�/3?�/W?�/T? �?(?�?L?�?p?�?�? �?�?�?SO>OwOO�O 6O�OZO�O�O�O_�O =_�Oa_�O_ _Z_�_ �_�_z_o�_'o�_$o ]o�_�oo�o@o�odo vo�o�o#G�ok �*��`�� ��1����*��� v���J�ӏn������ -�ȏQ��u����4� F�X����ޟ���;� ֟_���\���0���T� ݯx����������[� F�����>�ǿb�Ŀ ����!ϼ�E��i�� �(�b��Ϯ��ς�� ��/���,�e� ߉�$� ��H���l�~ߐ���+� �O���s���2�� ��h�������9�16 1�<���� 2������������� ��R��v�5 �Yk}�< �`����U �y/�&/��� /�/k/�/?/�/c/�/ �/�/"?�/F?�/j?? �?)?;?M?�?�?�?O �?0O�?TO�?QO�O%O �OIO�OmO�O�O�O�O �OP_;_t__�_3_�_ W_�_�_�_o�_:o�_ ^o�_ooWo�o�o�o wo �o$�o!Z�o ~�=�as� � ��D��h���� '���]�揁�
��� .�ɏۏ�'���s��� G�Пk������*�ş N��r����1�C�U� ���ۯ���8�ӯ\� ��Y���-���Q�ڿu� ����������X�C�|� Ϡ�;���_����ϕπ߹�B���f�L�^�7 1�i��%�_��� ����%���I���F� ���>���b���� �����E�0�i���� (���L��������� /��S�� L� ��l��� O�s�2�V hz�/ /9/�]/ ��//~/�/R/�/v/ �/�/#?�/�/�/?}? h?�?<?�?`?�?�?�? O�?CO�?gOO�O&O 8OJO�O�O�O	_�O-_ �OQ_�ON_�_"_�_F_ �_j_�_�_�_�_�_Mo 8oqoo�o0o�oTo�o �o�o�o7�o[�o T���t� �!���W��{�� ��:�Ï^�p������ �A�܏e� ���$��� ��Z��~����+�Ɵ ؟�$���p���D�ͯ h�񯌯�'�¯K���o�
���yߋ�8 1ז�@�R���
���.� 4�R��v��sϬ�G� ��k��Ϗ�߳����� �r�]ߖ�1ߺ�U��� y�����8���\��� ���-�?�y������� ��"���F���C�|�� ��;���_��������� ��B-f�%� I���,� P��I��� i��/�/L/� p//�///�/S/e/w/ �/?�/6?�/Z?�/~? ?{?�?O?�?s?�?�?  O�?�?�?OzOeO�O 9O�O]O�O�O�O_�O @_�Od_�O�_#_5_G_ �_�_�_o�_*o�_No �_Ko�oo�oCo�ogo �o�o�o�o�oJ5n 	�-�Q��� ��4��X���� Q�����֏q������ ���T��x����7��������MASK +1�û����~�XNO  ����MOTE  �3����i�_CFG� �p�����P?L_RANGl�g��t�POWER ��õݠ|�SM_�DRYPRG �%p�%m���TA�RT �ծ#�U?ME_PRO������_EXEC_�ENB  d�x�GSPDX�����;��TDB��Ϻ�RM޿ϸI_AIoRPUR�� p��B�<�ٛMT_�T�Рn��OBOT�_ISOLC1���8�����9�z�NA_ME p�n��ۙOB_ORD_�NUM ?ը�5�H844w g��b�w� ���w/(/�^/��/���PC_TIMEOUT��{ x�S232���1�4�γ L�TEACH PENDANPЅ��������l�j��Maintena�nce Cons�g��߾�"��f�?No Use���� ����0�B�T��h��NPO2�RҤ��z�e�CH_Lf[��p���	��~��!UD1:��z��R�VAIL���R����x�e�PA�CE1 2�p�
 �濫��{鋓Ć�����9˺�8�?�%���%��� 4IDu����� ��Y������) :!4�8�Uu�� ����/�) :/!/O/q���U/ ���/ ?�/?6?? K?m//�/�/�/c?�/ �/�/�?O2O	OOi? {?�?�?�?_O�?�?�O GO_._@_'_eOwO�O �O�O[_�O�O�_o�_ +_<o#oQos_�_�_�_ Wo�_�_�o�o8 Moo�o�o�o�o�o �o�D��4��I� k}���a��� 돽��0�B��+�X�2a�s�������W� ͏�����4�U�<�j�o�3~�������Ɵ t����<���Q�r�Y���o�4������ѯ 㯑��)�8�Y��n���vϤ�o�5��ʿܿ � Ϯ�$�F�U�v�9� �߬ߓ���o�6���� ������A�c�r��@V�������o�7�� ��(�:���^������s���������o�8 �!�3�E�W�{��� �����o��G �/ tm�
u d  /����� �/Nl -S-L/�/p�d� z��/ �/�/�/??&?/./ @.1:n?�;�?�/�/(? �?�?OO*O<O2?D? V?h?�?�O�O�?�?HO __&_8_J_\_ROdOpvO�O�O�_ ` @p��U]/o�O�IAakU�_Rodoj_ DjEowo�o�o�o�o�o %�o�o=A Se���	��� 3�E���+�]���a��o\
#o�o�_MO�DE  /
�S �/㏙_�ZA�oH�����	���㟐�CWORK_{AD�
����/R  /< 1����_INTVA�L�a�%�R_O�PTIONR� �%���V_DAT�A_GRP 2�,uX:D�@PП�� ̟�˩͏���1�� U�C�y�g�������ӿ ������	�?�-�O� u�cϙχϽϫ����� �����;�)�_�M߃� qߧߕ߷�������� %��I�7�Y�[�m�� ������������� E�3�i�W���{����� ��������/S Awe����P��$SAF_DO_PULS�Q�A���� CAN_T�IM��E}�R� ���Ƙ/qsy��֡��Yo�K�C  կ������l�//%/7/I/[/e��C�2�$K�)�d�$�!ѢIf) �P5��/�/�/���)�/� ��4�_ �R  T0�!?^?�p?�?�9T D���?�?�?�?�? OO $O6OHOZOlO~O�O�O��O�O�OU�s��'��O$_6_�I  }�T;�o���WQo�p�M
�t��Di��[=Z0 � ��o�[Q [SC�_�_�_�_o  o2oDoVohozo�o�o �o�o�o�o�o
. @Rdv���� �����*�<�N� `�r��������?�� я�����+�=�O� ��r%{�������ß՟������"�_���0 2�SwU�]n������� ��ȯگ����"�4� F�X�j�|�������Ŀ ֿ�����0�B�T� f�xϊϜϮ������� ����,�>ߩ�b�t� �ߘߪ߼�������� o�(�:�L�^�p��� ���#�Q�[����
� �.�@�R�d�v����� ����������' 9K]o���� ����#5G Yk}�������O�3�//1/ C/U/g/y/�/�/�/�/��/�/�/	??-?;:p�D?q?{6��d��j?@]	123�45678�Rh!B!����B��V��?�? OO)O;OMO_OqOwA ��O�O�O�O�O�O_ _*_<_N_`_r_�_�_ �_�_�]�O�_ oo$o 6oHoZolo~o�o�o�o �o�o�o�o�_�_D Vhz����� ��
��.�@�R�d� #��������Џ�� ��*�<�N�`�r��� ������y�ޟ��� &�8�J�\�n������� ��ȯگ����ϟ4� F�X�j�|�������Ŀ ֿ�����0�B�T� f�%��ϜϮ������� ����,�>�P�b�t� �ߘߪ߼�{������ �(�:�L�^�p��� ��������� ����0.�@�%���l�~�����Cz  B}\�   ��}2d4� ���d1
���  	�d22,�%7I�Xp���Z�� ����� %7I[m�� ������!/3/ E/W/i/{/�/�/�/�/ �/�/�/??/?A?S?e?w?�?�:Z������<�4��`�$SC�R_GRP 1��� �� ߐ ��� ���	 �1��2
BD [����� I�7GDO2O�kO�����hBD?E� DP�wC��GhK�ARC� Mate 12�0iC 6789�0��M-�@A }8��M2IA�A���
12345t�D;F�2  ����>U�1{F�1HC�1��AhAJ<ANY	�?R�_�_�_�_�_�\��H��0�T�7�2 o/O0oVoho7F/��Co�o?o�o����l0Q�o:DBǲ�Ɛr2tAA��A c @��YuA@�WpNj ?�wrH����DzAF@ F�`�r��o��� ��B�-�f�Q���}�Yq�r������ďքB��y�*��N�9�r� ]�o�����̟���۟ �&���CTOF�k������h�����qYq6'�裯7G@Ypݯ����W\HC+�3���AnpC�V��o�~ec��W���  y���������ո�\�¿ P�(�@%�7�I�v�b�SS��0�EL_DEFAU�LT  m�����u�HO�TSTR��d���M�IPOWERFL�  ������W�FDO�� �� �u�RVENT 1����`�� �L!DUM_E�IPL�(��j!?AF_INE��Fߞ��!FT�u��<ߙ�!o�� ������!RPC_OMAIN���غ�ߜ1���VIS��ٻ� �}�!TPp�P�Ut�/�dl���!
�PMON_PROXY��2�e��������+�f�a�!R?DM_SRVb�/�9gP���!RT���0�h����!
��M�,�,�i��E!R�LSYNCFl	�84�!ROS�߸�4��!
�CE��MTCOMd�2�k�)!	�OCONS*1�l�u!�WASR�C|�2�md�!N�USB�0�n�>/!STM��'/.�o�Y/��}/p�J/�\/�/�/�/�/��ICE_KL ?%�� (%SVC�PRG1�/::$52�:???)03b?g?)04��?�?)05�?�?)06�?�?)07OO)0
T$JOE<9ROWK&4�� O)1,?�O)1T?�O)1 |?�O)1�?_)1�?G_ )1�?o_)1O�_)1DO �_)1lO�_Q1�OoQ1 �O7oQ1�O_oQ1_�o Q15_�oQ1]_�oQ1�_ �oQ1�_'Q1�_OQ1 �_wy1%o�/	2)0? "0��I1�/��S� >�w�b�������я�� ������=�(�a�L� s���������ߟʟ� �'�9�$�]�H���l� ����ɯ��ۯ���#� �G�2�k�V������� ſ���Կ���1���C�g�Rϋ��*_DE�V ���MC:�Ƞ��~��GRP 2�����0bx 	_� 
 ,���� ߟ���7��[�B�T� ��xߵߜ�������� ��3�E�,�i�P��� ����z��������� A�S�:�w�^������� ��������+O ��D�<���� ��'9 ]D ��z����� /h5/G/./k/R/�/ v/�/�/�/�/�/?? ?C?*?g?y?`?�?�? �?�?*/�?�?O-OO QO8OuO�OnO�O�O�O �O�O_�O)__M___ F_�_�?x_�_p_�_�_ oo�_7oo[omoTo �oxo�o�o�o�o�o �oE�_i{b� �������� A�S�:�w�^������� я�����^+��O� a�H���l�������ߟ Ɵ����9� �]�D� ����z�������� ���5�G�.�k�R��� ����ſ���������C�*�<�yϟ�d ���	gϰϛ��Ͽ�0�����+�%�+�P������i��i� y߇�qߧߕ��߹��� ��=�"�e���O�=�s� a���������3� ��'��K�9�o�]�� �������������# G5k�����[ �W���C �j�3���� ���/]B/�/ u/c/�/�/�/�/�/�/ 5/?Y/�/M?;?q?_? �?�?�?�/�?�?�?�? �?OIO7OmO[O�O�? �O�?�O�O�O�O�O_ E_3_i_�O�_�OY_�_ �_�_�_�_�_oAo�_ ho�_1o�o�o�o�o�o �o�oIooo@os a�����!� E�9��I�o�]��� �����ޏ������ 5�#�E�k�Y���я�� ����ן���1�� A�g�����͟W����� �ӯ	���-�o�T�f� �?���������Ͽ �G�,�k���_�M�o� qσϹϧ�����C� ��7�%�[�I�k�m�� ������ߥ����3� !�W�E�g���ߴ��� ���������/��S� ��z���C���?����� ����+m�R�� �s����� E*i�]K�o ����/A� 5/#/Y/G/}/k/�/� �/�/�/�/�/�/1?? U?C?y?�/�?�/i?�? �?�?�?�?-OOQO�? xO�?AO�O�O�O�O�O �O�O)_kOP_�O_�_ q_�_�_�_�_�_1_W_ (og_o[oIoomo�o �o�o	o�o-o�o!�o 1WE{i��o� �����-�S� A�w�����g�я�� �����)�O���v� ��?�����͟���ߟ �W�<�N��'��o� ����ɯ���/��S� ݯG�5�W�Y�k����� ſ��+�����C� 1�S�U�gϝ�߿��� �������	�?�-�O� ���Ϝ���u��߽��� ����;�}�b��+� ��'���������� U�:�y��m�[���� ��������-�Q��� E3iW�{�� �)�A/ eS����y� u�//=/+/a/� �/�Q/�/�/�/�/�/ ??9?{/`?�/)?�? �?�?�?�?�?�?OS? 8Ow?OkOYO�O}O�O �O�OO?O_OO�OC_ 1_g_U_�_y_�_�O�_ _�_	o�_o?o-oco Qo�o�_�o�_wo�o�o �o;)_�o� �oO������ �7�y^��'���� ����ُǏ��?�$�6� ���W���{����� ՟���;�ş/��?� A�S���w����ԯ� �����+��;�=�O� ��ǯ���u�߿Ϳ� �'��7ύ�����ÿ ]Ϸϥ���������#� e�J߉��}�ߍ߳� ��������=�"�a��� U�C�y�g������ ���9���-��Q�?� u�c������������ ��)M;q�� ��a�]�� %I�p�9� ������!/c H/�/{/i/�/�/�/ �/�/�/;/ ?_/�/S? A?w?e?�?�?�??'? �?7?�?+OOOO=OsO aO�O�?�O�?�O�O�O _'__K_9_o_�O�_ �O__�_�_�_�_�_#o oGo�_no�_7o�o�o �o�o�o�o�oaoF �oyg���� �'�����?� u�c���������#� ����'�)�;�q�_� ��׏�������ݟ� �#�%�7�m�����ӟ ]�ǯ���ٯ���� u���l���E�����ÿ ���տ�M�2�q��� e���uϛωϿϭ��� %�
�I���=�+�a�O� qߗ߅߻�����!߫� ��9�'�]�K�m�� �ߺ��߃�������� 5�#�Y������I�k� E���������1s� X��!�y��� ��	K0o�c Q�u����# /G�;/)/_/M/�/ q/�/�/�//�/? ?7?%?[?I??�/�? �/o?�?k?�?O�?3O !OWO�?~O�?GO�O�O �O�O�O_�O/_qOV_ �O_�_w_�_�_�_�_ �_oI_.om_�_aoOo �oso�o�o�oo�o �o�o�o']K�o ��o����� �#�Y�G�}����� m�׏ŏ������ U���|���E�����ӟ ������]���T��� -���u�����ϯ��� 5��Y��M�߯]��� q�����˿��1��� %��I�7�Y��mϣ� ���	ϓ�����!�� E�3�U�{߽Ϣ���k� ����������A�� h�z�1�S�-����������[�@�����$SERV_MA_IL  �����e�OUTPUT�t���RV �2�	�  �� �(�O���i�SAV�E��g�TOP10� 2�� d ��;M_q�� �����% 7I[m��� ����/!/3/E/ W/i/{/�/�/�/�/�/��/�/??/?	�Y�P��f�FZN_C�FG �	����.��o1GR�P 2�y7�� ?,B   A�0.�D;� B�0��  B4.R�B21��HELL�r2�	���������7"O1K%RSR 1O2ODO}OhO�O�O�O �O�O�O�O_
_C_._�g_R_�_�_�^�  ��%�_�_�_(�R�\a. �_b�`ރ��R2. d�o�_�6HK 1��; o�o�o�o �o�o�o�o
3.@ R{v��������<OMM ���?2��2FTOV_�ENBt����HO�W_REG_UI�R�g�IMIOFW�DL��!��5A���*SYSTEM�*. V8.303�40 ł11/9�/2020 A� ���X�SN�PX_ASG_T�   0 $�ADDRESS � ��ZE�V�AR_NAM	��%$MULTIP�LY��PAR�AM�� � �$TIME����$�_ID�	$�NUM�D�T�CI{MP[�FRIFD�VERSION���G�TATU �$wDISK�NFOD��MODBUS_A�DR[�����POR�C�`�SSR��� x ��NG�LE��g�$DU�MMY7�SGL��TASK   &����T�������STMTT0�P�SEGT2�BWD��h��E��SVC�NT_GP�� �8 $PC�E�R_V�   �	$FB�Pm�ScPC��m�ΐVDX��R[�� �$DATA00��u���1��2��3���4��5��6��7���8��9��A��B���C��D��2���FP�� y���1Ω1۩U1�1��1�1�U1�1)�16�1C�U1P�1]�1j�1w��ҀI���2Ω2۩2��2��2�2�2��2)�26�2C�2�P�2]�2j�2w�3���3��3Ω3۩3��3��3�3�3��3)�36�3C�3�P�3]�3j�3w�4���4��4Ω4۩4��4��4�4�4��4)�46�4C�4�P�4]�4j�4w�5���5��5Ω5۩5��5��5�5�5��5)�56�5C�5�P�5]�5j�5w�6���6��6Ω6۩6��6��6�6�6��6)�66�6C�6�P�6]�6j�6w�7���7��7Ω7۩7��7��7�7�7��7)�76�7C�7�P�7]�7j�7w����S�PRM_U�PDӑ  9$4q� 
�����ӑؐ$TOR�QUE_CMD �  u�MOa_�SPEEjQ_C�URREo�nAX�I �mS�CAkRT��_Ut���̒YSLO� � �������������_�{�V7ALU�OP��$�#(F�ID_Ll��K%HIF*IN�$FILE_A��v$�$M�t��S}AR0  h^~� E_BLCK����"���(D_CPU �)��)��F#y/�$����_=�R 	 ߈ PWҐOT쁑)1LA#�SR� .3?184RUN_�FLGQ5-4U184W�ITX5v1-4v185H�2�D4�084̑TBC�2��
 � �$O�X0IGu �0_OFTM1D��42D�WTDCX0AZ��2aM���6�1�7TH��"C�DxGR.0A��ERVE�3?D�3r?D3O��0_AC@� X -$jALEN�3wD�3j@EL_RATI���$�W_�F#14jAc$2�GMO�!>�|�C��ERTIA�`o!�Iaj@�KDE�E���LACEM�CiC�CmV�@MA�p�F7UW7QTCV>\_QWTRQ^\UuZ����Ct��USt�J_$��q�M�TF�J2'��R�E�QUvA2�P`>�s�a�C@JKfVK�1'a�1'a`A`�J0<d+cJJ3cJJ;cAAL+ca`3c�a`[f4\e5C�PNA1�\�`Q[;P�L�@i_�E��3CF�� `^GROUP1 ����y�N�0CC�~�`REQUIR*B���EBUZ�fA�V$T�@2#qg@v��14 \�E�NABL	�$A�PPRpCL�
�$OPEN`xCLOSEozSE�y�E�
�1.� �u M��0<PPB�t_MGr!�pC��� �x��9P��wBRK�yNOL�D�vh�RTMO_��3���uJ"��P cdP3cP;cPcP�cP6P��S�b�Ց|�2�5� rđB�1���1��PATH��ӁɃӁ�Hσ�0�(p�W�SCA�Tr�ar�qINiBU�C�@��)�C��UM2�Y�@+@�P9�O!�EAT��0T�`@T�PA�YLOA�J2L�7R_AN�1��L�*0���������uR_?F2LSHR9DؑLO��(�ٗF��F�ACRL_�!&���"���4bH$ �$yH�rG�FLEXcsu�1J�6 PMr �?�?>OPO� c�iE :vO�FP ٧�O5aP�O�O�LF1�>�R��O�O�O�O_!_��E+_=_O_ a_s_�_�_�_�_Y�v� �W�Sdf����_�_ o$�jT2'W�X�`� eŴ��e'� �*o<o No``deme[ee�o�o�o�i�2J�d ���0�o�o� 8ATk�q�PELٰ}1=�jxJ(p#pJE �gCTR"�f�TNR�9�wHAND_V�B�c�0 �� M$��F2�v	D#�SW�!�3�v� $$M���yv�q����q�����>��A@R ���vQ!5��}A�| �zA�{A�@��{T� �zD�{D�P�G@0��ST�w���y��N�DYW0^p�v !�H���k@ϗ�ϗ�@��g������PX��a�j�s�|�������9 Ģ�� ��Ťข��qASYIM��^�p������_�0�.�A� +�-��K�]�o�����J��K�����˙x�_VI��	(�s V_UNIC.$P�בJeG"uG"�K$ �X$|&
��P�K�,��>��%�T�\��dà�0H+0Rr���!v�VrDI�sOp4�2� �c `�
O�I2AO�F�I1l��WW3o�~0�0ܰ�  � � ��M�E��@r2�"YT0PT���ڀ�1�`��du���8�1�9T���a $DU�MMY1`A$P�S_i�RF+�  tڀ�6XpFLA�`�YP��B�3$GLB_T��5*E�0�Vq�`��j�v1 XXMpw��ST±#p�SBR��M21_�VrT$SV_E�R��O� pC�CCL�D@pBAڰOL2� G�L EW� 4\�`�1$YQ�ZQ�!W�C`ԑ��As02�t��AU�E ��yN�@�$GIz�7}$�A �@�C�@� L�`V��}$F�EVNE+AR��Np�F]Y���TANCp���JO�G�A� ��?$JOINT
Ѻ`��"�@MSET��  WECU۱�S��'U��� �g�U��?�#pL?OCK_FO����0BGLVm�GL�hTEST_XM�cp�QEMP�Pr8+bBB�P$U���BF2�2#p�CQabh���PQarACE�`|Sr` $KAR�}M3TPDRA�@�d�QVEC��f�PkIUQaVaHE�POTOOL2��cV1�;RE�`IS3���b96s�f�ACH�P(p��aO��3�429��2�`ISr  @�$RAIL_BO�XE
��@ROB�O"d?��AHOW�WARO�Aq�0qROLM�2gu��
txrp��/pZ���O_F�Џ! �D�a� T�^�PR�`Oˢ!�R�*��Q�p�0�COU�R"XBMeYC���P$PIP#fN ���b/r�ax�Qa�p��?CORDED�P���q� ��OY0 #o D )@OBu� G��Pd�S��3(@S���I�SYSS�ADR8H�� �0TCH�SЛ ,0EN2�A��Q_T������P�VWVAu1% Ǥ �`�B5PR�EV_RT�$�EDIT�VSHWR��\F$����A%	 D�0��;���?$HEAD�� 4U���KE�A�0�CPSPDl�JM%Pp�L5b�R��44�&[�t���I,`SH�C��NE�`I��OTICK2�<M}���!��HNRA'� @]�����t�_GqP�&v��STY��qLODA�㖒��m�_( t 
 �GƅS%$�T=\@S>�!$=!2��1EF0rFP�SQU�`x%�B!TERC�0�Q���S��)  Ph@�׹���g��a�`1O�0�3t�IZDQE�1PRE��1!�̯��pPU�1�_DYObR��XS�PK6�AXIP��sVaUR�ڳI�Hp�~����_�`��ET��P( bl�O�FP�A�4 ss�`���SR��*lѠ�������� ���#��1��A� R�c�R�s�RŃ�d�~� ��dŢ������ː́C��|����!S�SC,@ + hƕ@DS��a�0SPLC0~�ATq��2��𐿒�2ADDRE�S�cB�SHIF��H`_2CHH�rz�IK@���TV�I72,��h���� 
+j
�rV�qA���'- \����O����<�C��򢵲����B<��TXSCWREEU�.	0k�TINA�CP��T��Q����� / T ���@����Ag@��^�p��^����RROL �wP��f���v��QUE���0 �� ��@S��A��RSM�T�U�NEX��6F�� S_�Cf�6V�i���6⒱C�RB��� 2-/��UE�1=2�B\��!�GMT� Li!�m�w@O�wBBL�_pW�0��2 ��O�O�ALE���GpTO�3RwIGH&BRD�D���CKGR�0NT�EX��OJWIDTHs1�u�"qA�a�%�I_�0H�� O3 8�!wP_T��ҭ�0R�@�RswH�2$� O�ѭ�4��I�GG U2 �R b�rqLUM�u���E#RV
��@� PaP���5{0�GEU�R&cF���Q)]�LIPM��E��C�)j@S�x�x�`w5u6u7u8Z���3��9P��6�a�QSv��4�USR�DO6 <���0UR���RFOC�aPP�RIαmp�!L T�RIP+qm�U)N$0547	Pt�$0���Yq��Hb���� q8�  �G \�aT�p1��ѣ"OS�1��&R���#�a�9��O�C�N�"�$�IaUU�:�/�/�U�N�#OFF!`��;[��3On0 ٰtW5�4:�@GUNw��P�0B_SUB8�2p@��SRT� �a<��vQ�p �ORpN�5RAU��4T�9䶇�1_���= |����OWN� T�$SRC���r�Dx!`CE�MPFI*�*ё�ESP-����� �e*B�&�b�!B�n��> `10WO8�rT�COP:1$��� _^@�b�A,�q�EWA�C?a�A�@�C�A�C �VC�CH�? �qC?36MFB1���Q�VC4�Y`��@x# %rT���XdP^Ȕ�spC�pRUDRkIV���_V��uT̐fpD�MY_UBY�ZTV��ħ�B��X�a�RP_�Sp�+��RL7�BMv$��DEY��cEX����EMU��1X7d[�USP�p�o��G��PAC3INΑ}�RGMAad�wbF3wb3wb���ARaE����a�r7S�wb�pA R�@G�PP�r�`5VR� �pB !d�_���2	�BN��RECcSWo`_A$pa�8c�O!��QA��1s�E�UB��� �q5VHKG�C��Iz���.p��zsEA���w�@� 1u5U�MRCV��D ��FOS�M� Cs�	p�rX3�c�rREF�� �v�v�q p7��p  �z��z��{;��vpA_@@�zq��{��S�/g�Sᡏ���8R��E �$�=�ߠ) �UӠOU��b��ZS @�e2�2��$��R� �ΐB��2Ѻ�Kq�SUL6s�C�@CO:�� 3D)`�NT�CZ���BY��e�!e�$�L��S���S�����!��JTǤFt +��ǱT� ��CACH+�LO����*`�����@ܣC_LI[MI��FR%�Tj��'���$HO� 6B��COMMpSB�O�0 ]�Ԉ�I؄h@V�P�b��_SZ3dn���6����12����[`��&����AaM]P�FAI&�Gvt���AD��BMRyEׄ9�_SIZ��PH�`��FASY�NBUF�FVRTaDk�w�I�aOL��SD_@3��W3P�'ETUc�QNp[��ECCU�hVEM�`��۲&�VIRC���VTP�pO���J�s�A�w�_DEL�A�cP�ƺ�KS��G��@9pCKLAS��3	ő_�F�ƀH$p"�S;��N��P/LEXEEI��B�/��4sFLK I  `]�^A��M���dwsP3S/�^@�bJ# ������#�#RS ORD@!��> 3 ނ)�UK��T\"����WwCb2V��g%L�`�Qۑ6D4��\*bUR4sp_R'�d��� ,a]��ծc�_od&� {g��`B*�T�'�'SCO��*�C� ad �"_f�"0�">�"K� �"Y�J_\_nZ��� �E\ AM�P�0 mPSMf%Mp"�%HADJT�/e���Bڒ� Np"q׬!L�IN]3q��XVR�h$O\���T_OV�R� �ZABCB�5P�bw�$��
O��ZIPg%Qp"DB�GLV�CL�R �ޘ�MPCF�5R � r ���$��QLNK�2
��-`|��S �|q����CM+CMi`C�CC�A�CtP_�  $J:4D��@Q J�V�4$0�tO΂UXW� ��UXE>a��E�[����	��u��TC ����r�YK�D"0 U�"���^IGHbcq�?(� �K��V g� vG��$B$���@1e�B�҉�&GRV�%�F� ���OVC �5�A7�w@�`���
VBI���D�T/RACEB�V�1�����PHER�P �W , �3I[�$SIM�A-Q� e#4P �e!V&��q�e!�m/!��%�៍/Kpb/t#_UN��@_+p&LC�д�% �%V M���ALIAS ?�e���%1�! ( he�!:?L? ^?p?�?�66?�?�?�? �?�?	OO-O?OQO�? uO�O�O�O�OhO�O�O __)_�OM___q_�_ ._�_�_�_�_�_�_o %o7oIo[ooo�o�o �o�oro�o�o!3 �oWi{�8�� �����/�A�S� e����������я|� ����+�֏<�a�s� ����B���͟ߟ�� ��'�9�K�]�o���� ����ɯۯ�����#� 5��Y�k�}�����L� ſ׿���ϸ�1�C� U�g�y�$ϝϯ����� ~���	��-�?���c� u߇ߙ߫�V������� ����;�M�_�q�� .���������� %�7�I���m������ ��`�������!�� EWi{&��� ���/AS �w����j� �//+/�O/a/s/ �/0/�/�/�/�/�/�/�?'?9?K?]?3�$�SMON_DEF�PRO �����1 �*SYSTE�M*p:RECAL�L ?}�9 ( �}d?�?�?�?OO0O �?UOgOyO�O �O�OBO�O�O�O	__ -_�OQ_c_u_�_�_�_ >_�_�_�_oo)o�_ Mo_oqo�o�o�o:o�o �o�o%�oI[ m��6��� ��!��E�W�i�{� ������D�Տ���� �/�S�e�w����� ��@�џ�����+� ��O�a�s�������<� ͯ߯���'���K� ]�o�������8�ɿۿ ����#϶�G�Y�k� }Ϗϡ�4��������� ��1���U�g�yߋ� �߯�B�������	�� -���Q�c�u���� >���������)��� M�_�q�������:��� ����%��I[ m��6��� �!�EWi{ ���D���/�///�*copy� mc:dioc�fgsv.io �md:=>172�.8.9.225?:142242/�/�/�/�4F"frs�:orderfi�l.dat vi�rt:\temp�\]/o/
??.?�,�&*.d�/�,�/�?��?�?�'
xyzrate 11 Q?@c?u?OO*O�%�7�?4 �?�?�O�O�O�$7�/�(mpba�ck�?xO__0_ [}.F#dbN0*�O��N�O�_�_�_�%2x��D:\O_�Pa_4 �y_
oo.o�!3�Ua �_�_nU�_�o�o�o�O �O^_�_
.A_�o�e_�o����"�$�SNPX_ASG 2 ����q�� P �0 '%R[1]@1.1��y?��#%�(�� L�/�A���e������� ܏��я����H�+� l�O�a�������؟�� ��ߟ�2��<�h�K� ��o���¯��̯��ۯ ����R�5�\���k� �������ſ���� <��1�r�U�|Ϩϋ� �ϯ�������8�� \�?�Qߒ�uߜ��߫� ������"��,�X�;� |�_�q�������� ����B�%�L�x�[� ������������� ,!bEl�{ ������( L/A�e��� ���/�/H/+/ l/O/a/�/�/�/�/�/ �/�/�/2??<?h?K? �?o?�?�?�?�?�?�? O�?ORO5O\O�OkO �O�O�O�O�O�O_�O <__1_r_U_|_�_�_ �_�_�_o�_o8oo \o?oQo�ouo�o�o�d��tPARAM ��u�q ��	��jP;tAp��h#t��pOFT�_KB_CFG � s�u�sOPI�N_SIM  �{vu��p�p�RVQSTP_DSB^~r��x�`�SR ay G� &(u�#��v�TOP_ON_ERR  "uJy?�_PTN �fr��A;�RIN�G_PRMI� ��`VCNT_GP� 2au&q�(px 	�̏p���ޏ���wVD��RP 1�i'p�y� R�d�v���������П �����*�<�N�`� ����������̯ޯ� ��&�M�J�\�n��� ������ȿڿ��� "�4�F�X�j�|ώϠ� ������������0� B�T�f�xߟߜ߮��� ��������,�>�e� b�t��������� ���+�(�:�L�^�p� ��������������  $6HZl~� ������  2DV}z��� ����
//C/@/ R/d/v/�/�/�/�/�/ �/	???*?<?N?`? r?�?�?�?�?�?�?�?�OO&O0�PRG_�COUNT?v�8r�NuRBENB��ME�MwCAt�O_UPD� 1�{T  
;Or�O�O�O__ (_:_c_^_p_�_�_�_ �_�_�_�_ oo;o6o HoZo�o~o�o�o�o�o �o�o 2[V hz������ �
�3�.�@�R�{�v� ����Ï��Џ��� �*�S�N�`�r����� �����ޟ��+�&� 8�J�s�n��������� ȯگ����"�K�F� X�j���������ۿֿ ���#��0�B�k�f��x�DL_INFO {1�E�@��	 ����������@���@���}?�¿���
���U�@�yߍ�� D����D��  6��´��ߞ�O@YSDEBSUG\@�@��d�I���SP_PASS�\EB?��LOGW ���C��9�ؘ�  ��A��UD1:\�<���_MPC�EH���AH�� �A~m�SAV �m�4�L��S�S�Vd�TEM_TI_ME 1	��@� 0��S�CKT1?SVGUNS�@]E�'�E�r�ASK_OPTION\@�E�A�A��_DI���xO��BC2_GRP 2
�I=���?@�  C�f��BCCFG ����� l�]`]`ߕ���� ���7"[F X�|����� �/3//W/B/{/f/ �/�/�/�/���,�/ �/"?4?�/?j?U?�? y?�?���?���0�? O �?$OOHO6OlOZO|O ~O�O�O�O�O�O_�O 2_ _B_h_V_�_z_�_ �_�_�_�_�_�_.oh � BoToro�o�oo�o �o�o�o�o&8 \J�n���� ���"��F�4�j� X�z�����ď���֏ �����0�f�T��� @o����ҟ���t�� �*�P�>�t�����f� �����ί���� (�^�L���p�����ʿ ��ڿ ��$��H�6� l�Z�|�~ϐ��ϴ��� ����2�D�V���z� hߊ߰ߞ��������� �
�@�.�d�R�t�v� �����������*� �:�`�N���r����� ����������&J  �bt���4� ���4FX& |j������ �//B/0/f/T/�/ x/�/�/�/�/�/?�/ ,??<?>?P?�?t?�? `�?�?�?OO�?:O (OJOpO^O�O�O�O�O �O�O _�O$__4_6_ H_~_l_�_�_�_�_�_ �_�_ ooDo2ohoVo �ozo�o�o�o�o�o
 �?"4Rdv�o� �������� <�*�`�N���r����� ��ޏ̏���&��J� 8�Z���n�����ȟ�� �ڟ�����F�4�j�  ������į֯T�����
�0��T�>�r���$TBCSG_G�RP 2>��  �r�� 
 ?�   ������ӿ������@-��Q�c�v�}����d0 ���?~r�	 HC�`��r���b�C�  B�����Ȣ�>�f�f�źƞ��������϶�\��H �h�BYLcφ�B$дh߀j߈ߎ߲߰����ތ��@�@��AƷ�f�y� D�V��������	�^�?333��2�	V3.00���	m2ia�	*T�L�q�c�"����r����� ���l���   ���B������u�J�2}���5���C�FG >���� ��
�D��o�o��
 G������� 5 YDV�z� �����/1// U/@/y/d/�/�/�/�/ �/�/�/????Q?�� ��\?n?�?*?�?�?�? �?�?O�?1OOUOgO yO�OFO�O�O�O�O�O 	_r�^�._:�>_@_R_ �_v_�_�_�_�_�_�_ o*ooNo<oro`o�o �o�o�o�o�o�o 8&\Jl��� ��������6� X�F�|�j�����ď�� ԏ����܏.�0�B� x�f�������ҟ���� ���*�,�>�t�b� ���������ί�� �:�(�^�L���p��� ����ܿʿ ��$�� H�6�X�~�(��ϨϺ� d����������D�2� h�Vߌߞ߰��߀��� ��
����@�R�d�� t���������� ����*�`�N���r� ������������& J8n\~�� ����"��: L
�|��� ����0/B/T// d/�/x/�/�/�/�/�/ ?�/,??P?>?`?�? t?�?�?�?�?�?�?O OOLO:OpO^O�O�O �O�O�O�O�O_ _6_ $_Z_H_j_l_~_�_. �_�_�_�_ oo0oVo Dozoho�o�o�o�o�o �o�o
@.Pv ��Tf���� ��<�*�L�r�`��� ������ޏ̏���� 8�&�\�J���n����� ��ڟȟ���"��F� X�op���o>�į�� �֯����B�0�f� x���H�Z������ҿ ��,�>���b�P�r� tφϼϪ�������� (��8�^�L߂�pߦ� ���߸�������$�� H�6�l�Z��~���� ����d����&����� D�V���z��������� ��
.��R@b dv����� �*N<^`r ������// $/J/8/n/\/�/�/�/ �/�/�/�/?�/4?"? X?F?|?�?8��?�?�? t?�?�?OO.O0OBO xOfO�O�O�O�O�O�O��O__>_(^  dPhS hV|_hR��$TBJOP_�GRP 20U��  K?�hV	�R�S�\��8P���p��Q�U � � � � �<�RhS @dP�R	 �C� ff  C�W�Q4b���<f9o >��ff\a<a=�Z�C�`���b�
&`H&`.g�o�gn�ѴW4e\e`b�o ?�a�d=�7LC�FnoBȂo#&`�`89u�o�c�33\uX�2h�P<��C\�vc@333@3a3|b}`�BL�w�HqDa�l�����u�Jh�p<X���B$�d��?�/��C*p��C����Z`y�x��k< ���q`?]`C�4.�ϏR�d��daG����{<g��L�]p@&b`yap�c�z{4ep�V��� �������ʟ���(� � �N��Z�����������ޯ��d�hV�0�4e	V3.0}0�Sm2ia�T�*Z��TcQh�s�� E�'E��i�FV#F"�wqF>��FZ�� Fv�RF��~MF���F����F��=F����F�ъF���3F���F��{G
G�dG�G�#
��D��E�'
EMKE����E�ɑE��ۘE��E����F��F���F��F�(��F5��F�B��FO��F�\��Fi��F�v��F��vF��u�<#�
<�t���@Ť� r_X�j�M�hTn�@��U�S��SESTPA�RSA�\X�P�SHR���ABLE 1��[��hS�ȃ� (�0cɞ�����gWToQ��	��
����T��hQ�����ȜC���RDI�ϬQ���� �2�D�Vվ�O ����������*���	S�ߪS ������� !�3�E�W�i�{����� ����������/ A�]�����̂	k�}� ���M�_�q߃ߕߧ����hNUM  V0U�Q�PpP� B�C���_CFG� P�a@�PIMEBF_TT��p��S���VERA�����R 1��[ 8e�hRdcP! 3P�  �  //$/6/H/Z/l/~/ �/�/�/�/�/�/�/?  ?2?{?V?h?�?�?�? �?�?�?�>��?O�:0OBOTO.OxO�OdO �O�O�O�O�O�O_,__P_b_�8�_�_�_�~_�_�_�_�_���_�K�@���MI__CHAN� �} mcDBGLV�����p`ETHERAD ?���`�n��?o�ox�o��p`ROUT�!p
!"t@|?SNMASK�h�>�a255.~uF��|��F���OOL?OFS_DI��GT� �iORQCT�RL p	��n��T�B�T�f�x� ��������ҏ���� �,�>�P�b�r�����������PE_DE�TAI�h�zPGL�_CONFIG �Qa��/�cell/$CID$/grp1��@3�E�W�i�{�1�	 ����ʯܯ� ���$� 6�H�Z�l�~������ ƿؿ�������2�D� V�h�zό�ϰ����� ����
ߙ�.�@�R�d� v߈��)߾���������}��N�`�r�������� ����)�;�M�_��� ������������l� %7I[m��� �����z! 3EWi���� �����///A/ S/e/w//�/�/�/�/ �/�/�/?+?=?O?a? s?�??�?�?�?�?�? O�?'O9OKO]OoO�O O�O�O�O�O�O�O_���User� View !�}�}1234567890B_T_f_x_�_`�_�T-`��_��(Y25Y�Ooo*o<oNo`o�_�_/R3�_�o�o��o�o�ogo)�^4 �obt������^5Q�(�:�L� ^�p�����^6�ʏ ܏� ��$���E��^7��~�������Ɵ؟7����^8m�2�D�V��h�z���럭��� �lCamera3Z)����(�:�L�*�E�v����� @_��ƿؿ�����  ̦�Y�^�pς� �Ϧϸ�_����� �Kπ$�6�H�Z�l�~ߥ�� ̦�i������� �� $���H�Z�l�ߐ�� ��������ߣ�Py�� 6�H�Z�l�~���7�� ����#��� 2D V���*������ �����"4F� j|����kͥ ��Y/ /2/D/V/h/ �/�/�/��/�/�/ 
??.?���l��/z? �?�?�?�?�?{/�?
O Og?@OROdOvO�O�O A?�� �1O�O�O
__ ._@_�?d_v_�_�O�_��_�_�_�_o�O�G9 �_GoYoko}o�o�oH_ �o�o�o�_�o1CPUgy�	Υ0�o �������o2� D�V��oz������� ԏ{�Ӡիx�-�?� Q�c�u���.�����ϟ ����)�;�M�� ΥA�䟙�����ϯ� 󯚟�)�;���_�q� ��������`��u��P� ��)�;�M�_���� �ϧ���������� %�̿޵���q߃ߕ� �߹���r�����^� 7�I�[�m���8�޵ �(�������%�7� ��[�m��������� ��������޵���I [m��J��� �6!3EWi  	�� ����//(/:/<L/^+   nv �/�/�/�/�/�/ ?? $?6?H?Z?l?~?�?�? �?�?�?�?�?O O2O DOVOhOzO�O�O�O�O �O�O�O
__._@_R_ d_v_�_�_�_�_�_b,�  
 (  }�( 	 �_ oo:o(o^oLo�opo �o�o�o�o�o �o$:�Z~* ̸i {� ����� �X5�G�Y��}� ������ŏ׏���� �f�C�U�g�y����� ���ӟ�,�	��-� ?�Q�c����������� �����)�;��� _�q���ʯ����˿ݿ ��H�%�7�Iϐ�m� ϑϣϵ���� ��� �!�h�E�W�i�{ߍ� ����������.��� /�A�S�e�߉��� ����������+�r� ��a�s���������� ����J�'9K�� o������ �X5GYk} ������0/ /1/C/U/g/��/�/ �/��/�/�/	??-? t/Q?c?u?�/�?�?�?��?�?�?:?p@  B"O4OFOCG `���)frh:\�tpgl\rob�ots\m20i�a\arc_ma�te_1�@c.xmlO�O�O�O�O�O�__(_:_L_XX�� X_}_�_�_�_�_�_�_ �_oo1oCoZ_Toyo �o�o�o�o�o�o�o	 -?VoPu�� �������)� ;�RL�q��������� ˏݏ���%�7�N� H�m��������ǟٟ ����!�3�J�D�i� {�������ïկ��� ��/�F�@�e�w��� ������ѿ������+�=�_H�1 �Oj@88�?�=�|�=�xϚϜϮ� �������0��<�f� P�rߜ߆ߨ��߼�����&��$TPGL�_OUTPUT �"H1H1 `�H�]�o��� ������������#� 5�G�Y�k�}�������@��������H�`����2345678901 2DVhz �>2����� �9K]o�}������ ��1/C/U/g/y/�/ #/�/�/�/�/�/	?�/ ???Q?c?u?�??1? �?�?�?�?OO�?%O MO_OqO�O�O-O�O�O �O�O__�O�OI_[_ m__�_�_;_�_�_�_ �_o!o�_/oWoio{o �o�o7oIo�o�o�o /�o=ew�� �E�����+�� �}[�a�s���������̍@b����h� ( 	  7�%�[�I��m����� ����ǟ���!��E� 3�i�W�y�����ï�� �կ�����/�e�S����^�w��� ѽ�����)�;� ��d�v�ϚϬϊ��� ��L���ߺ�(�N�,� >߄ߖ� ߺ���n��� ���&�8��D�n�� ^��������V�� "���F�X�6�|����� z�����x�����0 B��fx��� ��N`,�P b@����p �/�/:/��p/ �/$/�/�/�/�/�/X/ �/$?�/4?Z?8?J?�? �??�?�?z?�?O�? 2ODO�?POzOOjO�O �O�O�O�ObO_._�O R_d_B_�_�__�_�_ �_�_oo�_<oNoTb��$TPOFF_�LIM ���p�����qibN_�SVm`  ӄ�jP_MON M#���d�p�p�2ӅiaSTRTC�HK $��f�^��bVTCOMP�AT�hq�fVWV_AR %�mAx.�d �o Y�p��bia_DEF?PROG 3vb�%p��d_DIS�PLAYt`�n�rI�NST_MSK � �| �zIN�USER�tLC�K��{QUICK�MENA��tSCR�E`���rtpsc�t�{���4b��_��STzi�RACE_CFGW &�iAtx`�	bt
?�܈HN/L 2'�i}� �H{ nr4�F�X�j�|��������ĚޅITE�M 2( � ��%$123456�7890��  �=<�7�I�Q�  #!W�_�kp��� bs�ů)����_�� ����^���y�ݯ���� 5�%�7�I�c�m�翑� =�c�u�ٿ�����!� ��E����)ߍ�5߱� ����Yߧ������A� ��e�w�@��[��� ���ߧ��k���O�� s��E�W���c����� �}�'�����o�/ ������;S���� #�GY"}=� as����1 �U/'/���� ��_/	/�/�/�/Q/ ?u/�/�/?�/i?�? �??�?)?;?M?�?O �?COUO�?aO�?�?�O O�O7O�O	_mO_�O �Ol_�O�_�O�_�_�_ 3_�_W_i_{_�_�_Ko qo�o�_�ooo/o�o �oeo%7�oC�o�o ��o���O�Ps�N�ڄS�)�>S��  ϒS�� �����y
 ාݏď���UD�1:\���e�R_GRP 1*���� 	 @ �pY�k�U���y�����ӟ�������͑��2��V�A�?�   q���m�����ǯ��� ٯ�����E�3�i�W����{��������	�!����c�SCB ;2+o� \�Y� k�}Ϗϡϳ��������Y�V_CONFIG ,o�󁧏��M���OUTPUT� -o�>���Yߝ߯��������� 	��-�?�Q�c�u�;� �ߝ����������	� �-�?�Q�c�u���� ����������) ;M_q����� ���%7I [m����� ��/!/3/E/W/i/ {/��/�/�/�/�/�/ ??/?A?S?e?w?�/ �?�?�?�?�?�?OO +O=OOOaOsO�O�?�O �O�O�O�O__'_9_ K_]_o_�_�O�_�_�_ �_�_�_o#o5oGoYo ko}o�_�o�o�o�o�o �o1CUgy �'�9Ո����� �#�5�G�Y�k�}��� ���oŏ׏����� 1�C�U�g�y������� ��ӟ���	��-�?� Q�c�u���������ϯ ����)�;�M�_� q���������˿ݿ� ��%�7�I�[�m�� �ϣϴ���������� !�3�E�W�i�{ߍߟ� ������������/� A�S�e�w����� ��������+�=�O� a�s������������� ��'9K]o ��������� #5GYk}�����x��� ����/�3/E/ W/i/{/�/�/�/�/�/ �/�/?�/?A?S?e? w?�?�?�?�?�?�?�? OO*?=OOOaOsO�O �O�O�O�O�O�O__ &O9_K_]_o_�_�_�_ �_�_�_�_�_o"_5o GoYoko}o�o�o�o�o �o�o�o0oCU gy������ �	��,?�Q�c�u� ��������Ϗ��� �(�;�M�_�q����� ����˟ݟ���%� 6�I�[�m�������� ǯٯ����!�2�E� W�i�{�������ÿտ������,��$T�X_SCREEN� 1.����}ipn�l/`�gen.htm,�ϑϣϵ����$ Panel� setup��}�����0�B�T�f����ϝ߯������� ��n���?�Q�c�u� ����"�������� �)�������q����� ������B���f�% 7I[m������ ����t��E Wi{���: ��////A/�/��UALRM_MS�G ?L��Y� Z//��/�/�/�/�/ �/??$?B?H?y?l?�?�?�?u%SEV � �-�6s"E�CFG 0L��V�  /�@��  A#A   B�/�
 �?6�L� VOhOzO�O�O�O�O�O��O�O
_W�1GRPw 21	K 0/��	 @Ob_u I_�BBL_NOTE� 2	JT���l6�Q�8��@uRDEFPROz %�+ (%�? �_8��_o�_'ooKo 6oooZo�o�o�o�o�o��ok\INUSER�  �]P_�oI_�MENHIST �13	I  (�@ ��(/S�OFTPART/�GENLINK?�current=�menupage?,153,17�8����� r�}936�,�>�P�b� �ry���������ӏ� t�	��-�?�Q�c�� ��������ϟ�p�� �)�;�M�_�q� ��� ����˯ݯ�~��%� 7�I�[�m�}��Rlq� ����Ϳ߿���'� 9�K�]�oρ�ϥϷ� �������ώϠ�5�G� Y�k�}ߏ�߳����� ������1�C�U�g� y���,��������� 	����?�Q�c�u��� ������������ ),�M_q��� 6���%7 �[m���D ���/!/3/�W/ i/{/�/�/�/�/R/�/ �/??/?A?�/e?w? �?�?�?�?�����?O O+O=OOOR?sO�O�O �O�O�O\O�O__'_ 9_K_]_�O�_�_�_�_ �_�_j_�_o#o5oGo Yo�_}o�o�o�o�o�o �oxo1CUg �o�������? �?�-�?�Q�c�u�x ������Ϗ�󏂏�� )�;�M�_�q������ ��˟ݟ����%�7� I�[�m��� ���ǯ ٯ������3�E�W� i�{������ÿտ��������$UI�_PANEDAT�A 15����A�  	�}�d�vψϚ��Ͼ� )���Ϟ�R� �!�3�E�W�i��ύ� t߱��ߪ�������� /�A�(�e�L����\�� ��� ����� �2�D�V��� z��ό����������� 
q�.R9d� o������ *<#`���C� ��������P !/��E/W/i/{/�/�/ /�/�/�/�/�/?/? ?S?:?w?^?�?�?�? �?�?�?Oz�=OOO aOsO�O�O�?�O./�O �O__'_9_K_�Oo_ V_�_z_�_�_�_�_�_ o#o
oGo.oko}odo �oO&O�o�o�o 1�oUg�O��� ���L	��-�?� &�c�J����������� ��ڏ���;��o�o ~��������˟ݟ0� �t%�7�I�[�m�� 柣�����ٯ����� ��3��W�>�{���t� ����տ�Z�l��/� A�S�e�w�ʿ����� ��������+ߒ�O� 6�s�Zߗߩߐ��ߴ� �����'��K�]�D� ����Ϸ��������� �d�5�G���k�}��� ������,����� C*gy`�� ��������}�,ew����)S�W��/"/ 4/F/X/j/��/u/�/ �/�/�/�/?�/0?B? )?f?M?�?�?�?�?Q������$UI_P�OSTYPE  ���� �	 �?#O�2QU�ICKMEN  �KO&O�0RE�STORE 16���  '��?X��O�C�OX�m�O�O__'_ 9_�O]_o_�_�_�_H_ �_�_�_�_o�Oo0o Bo�_}o�o�o�o�oho �o�o1C�og y���Zo��� R�-�?�Q�c���� ������Ϗr���� )�;����Z�l�ޏ�� ��˟ݟ����%�7� I�[�m��������ǯ ٯ�����
�|�E�W� i�{���0���ÿտ� ��Ϯ�/�A�S�e�w��1GSCREA@?�FMu1sc��@u2��3��4���5��6��7��8<���2USER����2��T����ks���U4�5�6�7��8��0NDO_CFG 7K<;��0PDATE ����Non�e4B��_INFO� 18����RA0%}���Q�������� '�
�K�]�@��d�� ����������*L���OFFSET ;FM�Ë@ �b� t��������������� N�UL^�� �����&VO(�
L*�UFRA_ME  �d����RTOL_AB�RTp�ӈENB���GRP 1<��IRACz  A������	//�-/?&I/[/�@@U��iѠMSK  ���ӢNm%��%��/�_EV�N��$c�
6U�2�=I9hi��UEV�!td�:\event_�user\�/T0C�7Y?)�F�<L1S�PR1W7spot�weld�=!CA6�?�?�?�@�$!�/ h?&O[OGl�OJO8O �O�OnO�O�O�O_�O �O�Oe__�_4_F_|_ �_�_�_�_�_�_=o,o aooo�oBo�o�oxo��o�o'�o�j)6W�RK 2>@�88"�� y�� ��
��.�@��d� v�Q�������Џ⏽� ���<�N�)�_���~���$VCCMUҳ?\ݨ�MR�2�E8;<�"�	�j���~XC5G6 *����h֜ �5�i�A@�7 p? ȗ� ;[�e�Ȇ���ů�����^�9%A���ٯ*�� B���E��I�ѯ j�����]�����ֿ�� �����0χ��f�Q��cϜ�O����ϥ�ISIONTMOU?� ��ů�FU���U�(�� FR:\��\�u�A�?  ��� MC*�LOG�7�   UD1�*�EX[�E!' B@ ���Ҁo�r���o������d ��  =	 �1- n6  G-����Ҭ6,��<��1�=���:����n�P�TRAI�N����1�E!�Adt��͓G8; (�� :��S����������� -��1�?�Q�c�u���Й���T���_��REⲐH�����LEX�E��I8;�1-e���VMPHASE'  ���A����RTD_FILT�ER 2J8; ��R����� ��1C#�� t��������//��SHIFT6�"1K8=<���/p/3��O/u/�/�/ �/�/�/�/?�/?)? b?9?K?�?o?�?�?�?�	LIVE/S�NAP�3vsf�liv4�?�>�� SETU�0BmenuOO�?}O��OfB/%L����	|H{O�O��?�J� ��@-�AdB8
�����K�M�QR��S����	'-_�ME�0�ļ�/!M�OM �zWqW�AITDINEN�D����TOK C 噰\���_S�_�YTIM����
lG�_,m�_Ok�_/j��_/jo�XRELE�K_g���Q��֗Q_�ACT�0^h(q�X_N3� N��)r%�Ox_��rRDIS�0~�n�$XVR�B�O �$ZABCv͒1P�� ,��r��2g7ZIP�CQ����/�A�S��z�MPCF_G 1	R�J�0��w��a��MP�sS���<�q����8�F�?�  ���.d�������D��D���S���*���;B���f�~�n�ҟ�{���E�2�6��´$�6�>Ȇ�n� h�z�����ȫ�pt���T|��w�YLIN5DqU|�  �e� ,(  *)��:���&�c�J���n� ���Ͽ�#��s� (��!�^ϡ��ϔϦ� ���e�K� ���$��`y�Z�l��{��2V�+q đ������ �������٧�D����^�A���SPH�ERE 2W	�� �Ϛ�ߓ������<� O�*�<���`������ }��������I�[� 8��\CU��������pZZ�f � �f