��   ��A��*SYST�EM*��V8.3�0340 11�/9/2020 A   ���	�BIN_CF�G_T   X� 	$ENTRI�ES  $QW0FP?NG1FU1O2F2OPz �?CNETG  ��DNSS* �8 7 ABLE�D? $IFAC�E_NUM? $�DBG_LEVE�L�OM_NAM�E !� FT�P_CTRL.{ @� LOG_8	��CMO>$D�NLD_FILT�ER�SUBDI�RCAPDS4��HO��NT.� 4� H�9AD�DRTYP� A H� NGTHOG���z +LS/� D $ROB�OTIG BPEEyR�� MASK@�MRU~OMGD�EVK\SY�R�CM+ �;$�� ��QS�IZNTIM�$STATUS_��?MAILSE�RV�  $PLA�NT� <$LIN>�<$CLU��f�<$TOcP$C�C5&FR5&JE�C!�ENB �� ALAR�BF�TP�w#�V8 }S��$VAR)�M�ONt&��t&A7PPLt&PA� u%��s'POR �_|T!["ALERT5&�2URL }>�#ATTAC[0�ERR_THRO��#US29�38� CqH- �[4MAX?wWS_1�y1�MOD�z1I� �$y2 � (y1PW7D  ; LAu00v�NDq1TRY�6DELA�3z0��1ERSIS�!�2��RO�9CLK�8M8� ��0XML+ �#�SGFRM�#TC�P�OU�#PINoG_RE�5OP�!UF�#[A�C�"u%_B_AUZ�@��B�"�COU!�UMM�Y1�G2?�RD�M*� $DI%S�� J@Io/ }3 $ARP��)_IPFOW_x��F_IN�FAD� �HO�_� INFO��wTELs P~���� WOR~�1$ACCE� CLV��RF�!��ICE�0�QF  ��$AS  �S���Q��
��
�PqV�1m@�W�@����QI0AL`�_�Q'0 �X
�����P�����@Bb;eA��� #m��!�Q�zo���$ETH_?FLTR  �Y.`W �������!��k�� #m2�kRoSHAR� 1#i  Pvo,8dXG|?�c �������B� �f�)���M���q��� 䏧��ˏ,��P�� %���I���m�Ο��� ���(��L��p�3� ��W���{�ɯ�� կ6���Z��~�A�S� ��w�ؿ������ �� ��V��z�=Ϟ�a��� �ϻ��������@ߒg�z _L�11�mx/!1.{�0I���z�1���2551.�Ղ����@ey�2�ߒ��Ц߸�������3�ߒ�o��0�B�T���4p�������������5���_�� �2�D���6`����� ������������6A�MY�(MY��p��P� Q� 8�<r����� �%7 �Pg y�J�����	//-/���Ce w/b,Q/��/�/�/�/��}iRCon�nect: ir�c4//alerts�/9?K?]?o?5 �/�?�?�?�?�?�?�e0cP9a���? 0OBOTOfOxO�O�O�O@�O�O�O�O_�$�?3_�`("_[_�/_�_H�_�_����`a�i�R>j�U�Q�Qt)Y�eI DMZcan�$TCPIP[b��mi(`=aEL�`��e�Q��`H!�TB�o�r�j3_tpdb/ �m�vQ!KCL�o�kv_.��V!C�RT�o�oF`�d?!CONSG�j=�asmonL�d