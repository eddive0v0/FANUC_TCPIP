��  �A��*SYST�EM*��V8.3�0340 11�/9/2020 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  �  �ALRM_�RECOV� � � ALM"EN5B��&ON&! �MDG/ 0 �$DEBUG1PAI"dR$3AO� �TYPE �9!_�IF� ` �$ENABL@�$L� P d�#Uژ%Kx!MA�$iLI"�
� OG��f �%CAUSOd�!PPINFOE�Q/ �L A� �!�%/ H� �'�)EQU�IP 20N�AMr �72_O�VR�$VER�SI3 ��!COU�PLED� $�!PP_� CES( C p71s!Z3> ��! � $�SOFT�T_I�D{2TOTAL_�EQs $�0�0N�O�2U SPI_I�NDE]�5X{2S�CREEN_84no2SIGU0o?|�;�0PK_FI� �	$THKY�-GPANE�4 ~� DUMMY1d�TDd!_E4\A!R��!R�	 � �$TIT�!$I��N �Dd�Dd �DTs@�D5�F6�F7�F8�F9�G0�G�GZA��E�GrA�E�G1�G1
�G1�G1�G �@!�SBN_CF>"
� 8F CNV_J� ; �"�!_CMN�T�$FLAGyS]�CHEC��8 � ELLSET�UP � $�HOC0IO@� }%�SMACRO�ROREPR�X� D+`�0��R{�UHM�P�MN�B�! UT�OBACKU��0 �)DE7VIC�CTI:0�A� �0�#�/`B�S�$INTERVA�LO#ISP_UN9I�o`_DO^f7��iFR_F�0AI�NA���1+c�C�_WA�d'a�jOF�F__0N�DEL��hL� _aAqQbc?Yap.C?�Y`�A-E��#%sATB��d��AW{pT $DB� g"� =S�$MO�0B x!kq� \� ;VE~a$FN!�p�d�_�t�rdTM�P1_F�u2�w1�_~c�r~b MO<� �cE D [�mp�a���REV��BIL0�!XI�� �R  �� OD�PT�$NOnPM��I�b�/"_�� m�蘁H��0DpS �p E RD_E�L�cq$FSSB�n&$CHKBD_YS�r�aAG G�"$SLOT_�H�2��� Vt�%��x�3 +a_EDIm   � �"���PS�`84%$�EP�1�1$OP��0�2qc�_OK8ʂ� e0P_C� c��+dR�U �PLACI4!�Q���( �a�p9M� <0$D������0pB�UOgB,�IG�ALLOW� �(K�"82�0VAaR��@�2�sBL�0;OU7� ,yq�`�7��PS�`�0M_Ox]d���CF��7 X0GR`0�z�M]qNFLI�<���0UIRE��$ށwITCH�sAX�_N�PSs"CF_�LIM�t=�SPEED�!���P��p�PJdV���u�u�3z`�P6��ELBOF� �W��W�pH� ���3P�� FB ���1��r1���G� �� WARNM�`d܁�P����NST� CORz-PbFLTR۵/TRAT�PT `� $ACCQa�N �r�pI�o"���RT�P_S�r C�HG@I�Z�T(���1�IE�T�Y1�݀�� x pi#�Qʂ�HDRBQJ; #C��2��3��U4��5��6��7��U8��9s!k�M$��	3 @F TR�Q��$�V����C�FN�_U�pY�k�OpT <F �������#�I2q�LLEC7�>"MULTI�b�"��A!cj DET_��R  4F S�TY�"b�=*�)�2��o���pT �|� �&$L�>�+�0�P��u�!TO���E`�EXT�יၑ8B���"2����
�t k0F�RLƯ�r�q���� !D"��M��Qm� �蠋c0���"��G�1�ց�qM���P��! �����# L0	����P �pA��$JO�B,�ǰR�0�TRIG��$ d������ �� �K� l��弧�1qC`�0b% t���F� CNG0A�qBA� ��x��
�!v@��� ��z�0�P{`X�R·&ΰf��Pt�a�!��"J!�_)R��rCJ$�*(J)�D�%CHӽ��z@h�P�Z�@ '.�RO`�&�ס�IT�c�NOM_�`���S��pTE(�@�݉��P�ǭ��RA�0�2&"<�>�
$TFV w�MD3�T���`U(C1[�g�'�Hgb�s1q*E���\Ѕs�q�ŦgAŦsA�YNTt�q�P|pDEF�!)��G�PU8/@������AX��Ģ�ewTAI~cBUFņ��|psQ* � l�'�PI�)�P\7M[8Mh9� k6}F\7SIMQS)@�KEE�3PAT�Ѡ"�%"�"$#�"�L�64FIXsQ+ �ԭ�AdC_v�����23�CCIh��5PsCH�P�2ADD�6�,AE,AG,A!H�_�0�0_,@�foA)� ԀzFK� '�=$#�"�:�4E��, l���7@zpF�CE�C!F+H�S�EDIS�G�3�-z�P��MARG����r%�FAC
��rSLEW<���x;�,M��MCY.����pJB����
aC�W�v��U�W/ ����CHNS_EMP��$GE g݀!_} ����pP�|!TC9f��y#a���Nd�W#%I��r<��<�J�R�И�SEGFRfoPIOj�ST`�gLIN׃�cPV����!�$0�����b�'��b�B��1` +`��	��a	`�� �a�Pܠ��At��Py�Q�SIZ���ltKvT`VsE pz�y�aRS%� ��uc@Q{k�|�`�xZ``Ld�| `�vCRCɥ��!����t�`%�p9a˭9b��MINQ��9a7��q�D�YCk�Cz��le��50�Lp ��EV���Fˁ_leF��N����Q(۶�X%+4,��#{0|!VSCA�} AY��c1G"�2 �>�
/Ψ`_rU@��+�w][��i %�7�2�;QR��3� @�ߒ߱���5ġR��HANC��$LG����*1$�0ND,�סAR�0NK�a0�q��acm�ME�1���n�A0h�RA��m�A�Z����X%O`�F�CT���7`�vS\�P
ADI�O� ��u��pWP �����Ā��Gv�BM�P�d�p�D&ah�AE�Sf@̓�W_P�B�ASk�s��4 � �I�T�CS�X@�w�5��	$��1�T��?sC�b�Ny`�aBP_HE�IGH71��WIDl�0�aVT�AC���u�!AQP0� �\�E�XP+�L�@��CU��0MMENU��6n��TIT�1	��%��aǱA1ERR9L���7 \���q��OR�D��_IDzG��QUN_Od�>�P$SYS���4��ő�Iϡ	�EV�G#�a��BPXWO�����8��$SK��*2 ��T(�TR�L��9 �� AC�`�u䈠IND� DIJ�4 _Z�*1KԬ*�W�PL�A�RWA.�tТSD�A�ת!��r@Y�UMMY9�ª�10���¾���:	�A1PR�q; 
��POSr��g; ��[$S$�q�PL��<��H�S@��=�'�C��>4�'�ENE�@T�{�?S�S��RE�COR.�@H ��O�@;$L��<$��62����`�_q�b��_D9�W0R	Ox@�aT[���b��.�F��������PA�c���bETURN,�V�MR��U� ��;CR��EWM�bmA�GNAL� 72$L�A�e��=$P��>$P٠= ?y�A<�C���@�DO�`����:���GO_AW ��M�O�a)�o���CS�S_CNSTCY�@A L� ^�C`'� ID[^�2
2
N��O���ـ}I�� B PNPfRB^rzCPI{POvI_BY�R�}�T�r��HND=G.�C H�DQ�kSP�s*�SBLI�O�F��0��L�S�D��0N0�	FB��FE��Ch��жE�DO&a-sO�MC`{�4(�C�rH��WFPBw�Z��SLA�P�F�bIN� �N3����G� $$���P]��v�� v�ޕ���!o�"�#ID�&L�&W��";$NTV*3"V9E 4��SKI��aHs�3�'2�b&aJ�x&aM�mdSAFE,d��'_SV��EXC�LU7ѻ���ON	L`�#YcL���4�ΤI_V8���PP+LYy�R��H[0'�3_M@�NPVR'FY_S�2MS�!O@��k6�1�~32�#Ot !5LS�E��#35�£1�`%�P��$��t5�%�g Hy��TA2МDP�� ҄S�G� I � 
$CURB�_�
� B�������#H��3F��UNM��DZD@���l�{IxA�X�J�F�EF��IM�J @�F]Bk��pOTb�k�ԋѭ5��h�P�и@M� NI��!K��
RwPA!(T�DAY��LOAD�j��R�ӵ2 �E�F/�XILy�Ĉq}�OhPe�D�_RwTRQ�QM DF����P�r�S`�ThU 2L�`���Qkp�P���Q�QN 0�A��QA�t�R���DUtb���"�CAB�a�O�B�NS�QW`ID�`PW���U/q� �VjV_�P�P����DIAG�1�aP�� 1$Vb�HuT�l��u�t� �j���rR�p�DQ�tVE��Y@SW�ad�p7`q�d�U�PM�p�QOH�Uf�QPP�`�sIR���rB��Fb�S��q��q �@3r��-x ��-uj�#e�PO��P���uR7QDWuMS���u�A�u�b�tLIFAEZ��C�p���rN�q �r�uxA�s�rI�xB�Cp���NC�Y���r�FLAW�y@O�V���vHE'ArSOUPPO2���rbS�_E�)E�_Xf�(h���s�Zp�Wp�p�`s���xA���XZ������qY2ˈC
�T������eN됕exAJJ� v_��q���/���Q `[ CA�CHE��3�SIZ��v*��"j�N� UFFIo� �p����Ե3��6����Mܞ���R 8�@KE�YIMAG*�TM��ᄣ��D��q�>��OCVIE�`�'S ���Ll$@)#?� 	��%����T�P�ST� !��`!��@!�VP!�|�0!�EMAILy��1Q��� _FAU�L��U� �9��C�OUz ��T��|aV�< $��zS��PC`IT�#BUF@F�)!F�Oy�o�D�	B��nC($�������SAV�Ţ�`� ��`���|FP
�z���d� _���"P_�#OT�����P[0���� B��AX��-�I����Wc7�_G�s��YSN_$q'�W�RDuTY��#rMb�T��F+�fP^@D�&�X������g�C_��&�K��8�4B�3��R��2�q��D�SP���PCy�I�M�pÖ��#�Æ`U`M�:���K0d�IPm#0�q	�o�TH��=�c�mPT��p�HSD=Im�ABSCz$��o�V� �Я�&�`��QNV�!GO�&ԑ�$mƸ�F�aаdR�����,�SCxbk(�M�ER4�FBCM�P3�ET�1�Y6��FUX�DU���\���%2CDf���z��u��R_NOAU]T�  Z�P4 ��"U�IUPS�CJ	@�C�1ϱב�㍰��[H *�L t�3���֚@ �0�#�����A��VQ���1�扑��7��8B��9���p���1��U1��1��1��1��U1��1��1 �2��2���2��2��2���2��2��2��2* �3�3��3���3��2����3��3���3 �4�_�X9T�aQ\ <2`�� �I簉���3刡�FDRxd]T��V�0���r��r�REM�`F��rO�VMI�>AGTR�OVGDT�gMXvING�fua'IND��r
��а$DG��:sp���u�aD�VpRI�V���rGEAR�I�IO�eK7�tN �%(hQ�x0h `��sZ_MCMÀ�qv;�UR��^ ,�b1?���� ?� .�a?�!E�0�!!����_P}p5P���`RI�դ$��aUP2_ ` VPģTD���3�#�?@�!�'�%�ŢBACܲa T�ŢڠZ�A);@OG.5%�C8T����IFIq�0��x�:pC5PTV����FMR2
b� �3LI ��3#/5/G/^|���u7_���R_��A�԰`M�/-D�GCLFuDGDMY_HLD�!�5�vP��tz3�c�P�9? T�FS]��d P2`�B�0��а$EX_�A�H�A�1kPl���@3[5�V�G:�
e �����SW�O�vD�EBUG4WR�eG�R� �U��BKUv��O1a� pPO�P�YoP��BUoP�MS�0OO���QS�M�0E���� _?E f �`����TERM�Ug<�UH��ORIe0�Qyh�U��SM_80�Ţ�Pi�W�TArij�U���UP㒟k� -���f$�Ua`g$SEyGfjx@ELTOV��$USE��NFI"��bn �q+�d>]dh$UFR02�`��a���	@OT�g�U�TA ��cNST`PAT��?��bOPTHJ ���E�8:��АbART+��ep|�+�V��aREL<z9�SHFT�a q..x_SHI�M^���"f $`�xj)A�0�OVR��ǲSHI�_p&DU4� %�AY#LO��AֱI�ѻ#p qk�%�k�ERV�� �q�yz��g`<r40_0&���_0RC�!9��ASYM	�9��aWJ�g��E�#*qV���aUz�`ֱ.u|����DuP���pYѪvOeR`M�3Z�GR�Q1Tl�oR�V�`�`A8��B��m �>�b6]71TOC�a�QT!k�OPZ2���}���303OYߠR%EM�Rm�9�Oѐ$�reT�R�e��h�|Fq/4e$PWR�3IM���rR_C�#t�VIS`sb�UD��#fsSVW�B��b ;n� $H.56�__ADDR�H�QAGr2�'� �
�R��\~�o H�@S�� Q�4_���_���_���cSE�A�HS���MN�Ap �T���_����OL����v���ּPAC�RO���aS�ND_�C����qٔZ�RO�UP���_X���@��1��25���?� 4 ?�<@���?���?�l��2AC�IO�ӂW�D:���J���1Sgq $� ;�_D� x�PM���PRM_.�}^�HTTP_��HQar (�OBcJE��"�/4$��LE�c��s � ���AB_��T�SS�S� �D�BGLV��KRL~ÙHITCOU�[BG��LOF�R�TEM�ī�xe�a7�f�SSQ ��JQUERY_FLA��G�HW��aQatZ����F�PUR�IO�h����u�у��ѿ� �IOLN�2u��
@C���$SL�2$INoPUT_�1$��bi�P m�D�SL��Qav��gߢԝ�=�s��=��QIO�F_AuS�Bw%0$L:0'�:1�q��U`|p�aaTժ�_��pHY�p ���^���UOP�Ex `��>������hᣐP�Ã�^�Ђ���x�� UJ�	y � � N�E�wJOG�g��D�IS�3J7���J8��7!PI�a���7_LAB�a3������APHI� �Q��9�D�@J7Jx�� �@_KEY� �K�LM�ONQaz� $X�R����WATC�H_� �s98��EL�D.5y� n�E{ ���aV�(���CT�R@s����%R� LG�|���DS?LG_SIZM�� `&�@%��%FD0I$;�Q2#�P= /" _�+��@���@�R ��P��S���� �ťV" ZIPDIU�r��N��3R}J���@P�A��]�d0�U�-�L6,DAUREA��/��h^GH0��!��B�OO2~� C��ӐIT�Ü>@���REC�SCRN�����D����'�MARG�2Ҡ�����N�H"����S3���W����A��JGMG'MgNCH����FNd�J&Kp'PRGn)UqF|(�p|(FWD|(�HL�)STP|*V`|(e0|(�|(RS�)H�+��C�t�#y���1P#'G9U籐$"' �r0&���"G`)WpCPO�7�*��#M07gFOCwP(EX�חTUIn%I�  # �2,#C8#Cl p!�p@��v3@���p�NࡎsANA�҉b�pV�AI��CLEA�R�vDCS_HIP\T�Bu��BO�HO�G�SI�G�HS�H(I�GN; ��Mm!��T�٤�@DE�(4LL�\�C���BU�PR`j���pT4B$1#EM������rR
Qa����pW��Ρ�4�OS1zU2zU3�zQYT�AR`� �����΁�esԲs�IKDX�P�r��O�PX��a�VST?�Ri�Y��a �$EfCkW��&f9fq
�U��V�� L�� �_�#�|p��U���ו�E��֕YU�_ � �� .������c �MC �{ ���CLDP?�>J�TRQLI�[�8���i�dFLG���`���srAD��w��LqDutuORG�� !21r��vyxu��t���dд� ���t"5�du� PT�`��bp��t�vRCLMC��t}��y����MI������ d)�QR�Q����DSTB�P��P [��h�A�X�bi�k���EXC+ESy� ;�M��U�%�O��d0;��jV��Z�]�_AW��\��������`KB�� \�����$MB���LI�I�REQoUIRE�cMON�<
�a�DEBU��;�uL�`MA� ڰ� ᛐ����q;�ND>S��'��fړDC�2:IN��7RSM�����@Np���F3��PST�� � 4}�LO�C�VRI���UEX�\�ANG�RY�;�O�DAQA�K�$t�1RBMF��]����Y�b0�eǥC�SkUP�e��FXS��IGG� � ����b�wÓc:6�d���%c�?��?�x.���DATACW�k�E��E�����Nn"R� t��MD��I�)���@��-����Hp��ᥴX�!�ANSW!��`Q�1��D��)$~��� n��� ÀCU; aV� px���LOj"�����5�W�3�E���U�M�;�RR2>B��� (E�N�A�q d$CA�LIa��GvA��2�9�RIN� ��<$R��SW0���)��ABC��D_J2�SEu�Y���_J3:��
��1SP���Y�P���3�"��
Y�J�J�CZ՞r��O!QIM��(�CS�KPz��1oC��Jq(�Q�ܺՠպհ׎e�_AZ�rV���E�LQU��OCMP0s�)����RT���G�1���5��P1��9�f�G�ZE�SMG00}��Օ`ER���Å�PA �S(���D�I�)�JG�`SC�L����VEL�aIqN�b@��_BL�@Y����Z�J���������YPIN�ACcR���	"x��f`_u�!�<���<�b܂�F���YPDH��t;����iP$V����'A$d�b�ȏP`��qy�B��H �$BEL��||�_ACCE��� �����IRCi_����ppNT�Q��S$PS���bL��� (s�	1<w@
PATH��_D��_3..���_wQ �� ��rb�CC ���_MG !$DD���`�FWE�~���������DE�P�PABN6ROTSPEE�{Q�`��{QDEFb���?$USE_��BC%P��C�0BCY��Z�q s�YNA�A�p}yм�}MOU�NGRR� O��Q�INC�m���h�x���i�ENCS���d�Y�&��f�# IN��RI.%���NT�����NT23_Ux��`�A#LOWL�AA~0��`�a&Da0@Y�C���`���C,��(&MOS�@�MO��ǀ�wPERCH[  ~#OV�� �' �Q�#F�d"&�F��
�gm �@w�A. 5L ADw��v�)%�d*_6�z&TRK���QAY I�3쁏1.�5�3n�p�����PMOM B�h��sp"�W����0�3azR��DUЋ�S_BCKLSH_C.!E��&� ��-�?D�JJ���CLALBP'"�q�0܀|E�CHK�`�US�RTYJ�N����T:Seqr}�_c�$_UM����IC�C����C(LMT�_Lwp� T̱WE]&P[P !U,�5A�+0gT8PC�!8H�`|��2�EC�p�bXT���CN_��N���V�SF���)Vg�a	'�|�Q.
e�XCAT�NSH������eq�
A
&F�/F�Z� P�A�D�_P�E�3_ �`���6� �a�3�d�E�JG�p���cO OG|�W��TORQUY /Ւ#�9� ?��"��� r_W�5�4C��<tP��;u��;uIC{IQ{I��F��.qaҐxp�� VC��0b�Z��r�1�~���s��uJRaK�|�r�v�DB���M���M�_DL��:2GRVBt;���;����H_L��b �i�COSv��v�LN�p�������d�@��mq׊Ō�q�Z����&�MY�����T�H��6�THET0j%NK23��`��㶣�CBe�CB��C��AS���mt���󌘑e�SB��p�GTS��(C�m�=���cM��ԃ$DU��@C7����� ���Q�F�s�$NE��ؠI@���C)���T�AX������h�s�s�LPHv�_�9%_�S�ңŅ ңԅ_��������EV��V����VʪUV׫V�V�V�V�V�H��E�²P��?aٸ׫H�H�UH�H�H�O���O��ONɹ�OʪO�׫O�O�O�O
�O�F_�����Ņ��Ė�SPBALAgNCEQԃQLE͐H_X�SP�9��ņ9�ԆPFULC�=�d�L�d�ԅ&�1���UTO_�@�eTg1T2����2N�A ��?�Ԗ��1f�D�5���1TP0O����,p�INSEG��!R�EV�փ "!DIF�y5K�1�0��1��l0OB&�lAE��72�p?�A$�LCHW3AR��AB�a�5?$MECH��%�X���FAX�1PJTp��z���З 
��q�%ROB� C�R(2��R���MSK_���� WP ��_WR���r0�?{41	b4 2`0�1#JD0���IN���MTCOM_�C�p��  �� 8�$NOR�E$#���t����� 4�0GRr��F�LA�$XYZ�_DA��nC DE�BU�� ��t��u 0�$uCOD[AG ���2���0�$BUFIND�X2 ��MOR#�� H-��0����FB �0�JD$���c�QVPTAA�+�2G6� �� $SIMU�L�` 13�3O�BJE;ТADJ�US�� AY_It�A	8D�OUT�`����0�_FI�=@T+p4 ��X�3p3�A�5DNrFRI(CXT8E�RO�` E3q[0��OPWO�p'�}, SYSBUq�( $SOP��A�U�3�PRUN,v��PAC�D��℟0_� NR�X�A�B��PP� IMAG�[A-�G�P�IM�Y"$IN,��!#RGOVRDM�� ��P   #`W�L_`��an%�B�PRB5P�X�`QMC_EDT/ �� PPNq�M�"<OQ@MY19NQ+ �M!SL;�'� x $OVSL��wSDI{DEX�S��&�SP1�"V3p�%N 1q�0378�"xA*M!_SETp'� @�0K2��AASRI�� 
^6_��j7�1v1+ 5� �P� �<T���`A�TUS@$TR�CI�H%�3BTM$�7�1I��$4NQ�3\� '� D-�E��"�2z�Ev��1!0l@�1EXE�0�A�!B*B�4S3�Z0.��03UP��9A$Y�' XNN�7�q�$�q�9� �PG���? $SUB�1����1�1�3JMPWAeI,`P	3�ELOP����$RCV?FAIL_CH��AR-���Q�P�Tx�U�R_PL�3�DBTB�a�R�B3WDV��UM�`T�IG�( ��4`TNL(`TjRRm���`$
p	1XQ� E�S�T|�R�ADEFSP�� � L-���Pq_�P��SUNI#��7�PmAR1@��3�_L�P�1* �@w�&�����`�� "<0��)�:T"NU�KETb(p���`P^R&� �h� ARSIZE����1��naS� O�R�3FORMAT���TTCO� ja�EeM���d�SUX��2�1PLIOR&��  $��P_�SWIu��!�fL�LB&�� g$BA�`1�ON9A�KPAM�0=y��BGAJ5���2r68v>��_KNOW8cNrA�U9AߐDx� �P9DC�ryPAY�[�t���y��wZ�sL��1��U!PLCL_~$� ! �sP,qv�tb"�vF�y�CRPO�z�2�tE	S���wR4��w�t/BASE$�J��W�S_J�qK�mA���fBu��r�q_T0��MAX4P�`AL?_ � $�Qh �1q�!��C[�D�sE�fr�J3����� =T� PDCK� ��>T"CO_J3����`��
�hr���� ����C_YQ�  � ��� �D_1�z2�tD���n�^���m�^|TIA4��5��6[�MOMS ��ȓе�ȓ��B�@ADਓ억��PUB�{R͔������e#��` I$PI�$�QM�=q�wk� B1�yk���������iqRM�q�!Ħ~AĦ�A�
��9d5SPEED�G�b��E�T ��T�EP-�C��pQ+�Q�ESAM(ЀE�����Ep{� m�$�� k� ~@Ƕ�P_�ֹm�k�v {��ŵ��,H��ǳIN̚�c��1����B�W�.�W�w�GA�MM��1��$G#ET9" �D;�u=
��LIBRcA�R]I��$HIb@_=!H�0k���Eh ��A����LW��4�+��@X��7���wP��CEUxv�[ �0 �I_b�xu��L��������ȓu��ٞ� ��$Ј 1U���I�0R��D\�0��kAT��LEf�=qЊ1M�7�ୄPMS�WFLTM��SCRsH7�����!��~Bv�dSV&�P� �A �����#S_SaAqs$��eCNO;�C�1fB<�����K�� ���S�C���hrǥ��m�D� a���� ��� в����U!C���X�����s �dMJ�߰ � ��YL(i�K���^SJ�| v!6O�K���BK��- ��OW�� �9���M$P���p����Dc�"��1�~B�`M��T2� �� $-�$$W� �%ANG"�q�  ����!��5P�&��o����c�#��X`O"���Zz�`�@n� �y�OM��+�(�:�L�^�p����CON@�U �c;�_�B� |ၰ��ș @&��@&�࡚m'X&��.��� B�$"�⥴`X$$Pma��PM0QU�� �� 8#`QCOU����QTHYPHO�/� HYS�`ES�-r� UE� ��S`O��d�   $P��@�Ŋ2UN�0br�@O��  � P�p�45�E��C�RROGSRA�1A2DO4�45IT�Ё1F0IN;FO�� %0g;��1A�aOI�2�{ (�SLEQ�� �1��0k6E1S�НD�� 4#`ENA�B"20PTION��C�T̢/G�TCGC]FA� @#`J$P���<2���RdH�0OBG�2S_ED��@  � �{K��q�3��E)�NU��G�HAUT�ECOPY�qI0�L����M��N�@�K��PR�UT �BNV@O�U�b$G92DT�aRGADJ��fbbX_ �R$`(pV�pVWnXPnX[��pV�`Pz�N��_CkYC"ZSNSE9�$ ��LGO����NYQ_FREQ�0�Wb��a�d23L��p�b�PnQÓb��5CcRE���#��IF���s3NA��%?d_}G��STATU' <��*7MAIL��YsyIN��$LAST�a����TELEMA�� �GFEASIA����H �b�1 ���f;B����I�0����R=q�!� R�rAB$+A��Ex0�V�a7vW�Cy��1�U8�I0�p�d�lvRMS_TRs��@��sr7��z��aktB�R��/ 	�b 2� =�_+��ve��w�r�� �fe��c�G�D�OUa3;�NHC�RP�R	 @��2GRIyD�1+CBARS��sTYC�ROTO�R��³�&0_[d!�P䂂B�OxD� �s �0�PORa3���[���SRV_`),˄ÆDI�T^�䁠�������4��5*��6��7��8��Q�F��A�#0$VALURs���d�q_�>D�� E���u1��aa��=@AN��㉒qaR�@a��T�OTAL��1��P�W�SIJ���REG#EN����#XxxI30e%!��� TR^s0����_S��^���CV nQ�D��B8rE�cN���!��42�@ÓV_H�k�DA�~���S_�Y
�rfS��AR��2� <RIG�_SE�ch�Â�e_�80��C_v�`�EN�HANC�!� �p�qEqb�ý�I#NT��� F.3�MASK��ipOVR�#P� N��`a
�_�*6^�M��B[��f�8��SLG����� \ ��eH �d��Sq�dDE⁁U��*7Ő�%��U��Q�TEj  �G (7��҆�J϶<�"cIL_M!d��P㈠�TQ� �Ë1�rpj�eV��C��P�_��op��M��V1V��V1��2�2��U3�3��4�4�� �ᄠ�������s��;IN��VIB� �Ĩ�����2��2��3*��3��4��4�ؾ� ��#"�������%���،ՠՌ�PLv`TOR� ��INb������  �p��MC�_F� 	���LP����B�ڐM�IB����#� 1 �)����KEEP_HNADD��!��<p��	C�_`�䂁��H ��O�!��P������\G���REM���쑥�;�R�W�U[de���HPWD  ���SBMo���G��1�2�� H COLLABu��a�������ؑEb�0I�T���0��� �,� FLbq$�SYN��M�C���d�UP_DL�Y��#2DELAhJ �nbY� AD�}�!QSKIP�'� Ļ�60ODD���t P_60_2�g0 ^ ����		Q�	�� �	%��
2��
?��
L��
Y��
9�Q�J2�R�P��CX]pT�SY��X]P��Y8�1���PRDC��b� ��@ReCg�R�4ae��"d��RGEpr@sl�:�FLG�!�Pa�SW�I��SP9C�3�QUM_Yt�_2TH2N&�# ~L 1� ��EF�@11�!� �l�����C��AT4�ET1��7s"k0o4�j!�@Y�j!<3\�HO�ME�"�P<$2D"рJ/\/n/�/�/�/�'3D"��/�/�/�/?!?
�'4D"�D?V?h?z?(�?�?�'5D"��?�?��?�?	OO�'6D"Հ>OPObOtO�O�O�'7D"ֻO�O�O�O__
�'8D"�8_J_\_n_H�_�_�%S��1�9 �q=#$���< T�-E��ٷ��LbLݖJcIOq�jiI�P���;!POWE��G� 4` wGb�ה ��b$D;SB�GNABqՔ�E C) ��� �RSw232Pe� ���U�P�ICEU�Qrt�E3 ��PARsITáՑOPB��޵�FLOW�TR``�c�3���CU+pM��UXTn���U��ERFACtC�UvѐFbSCH�q'� t����_p�f�$����OM۠�9�A�T>���UP%D�A#�`T+`҃�*�� �x�s!��FqA������RSPqp�Q��� !�X$USA ���Y�EXmpIO6��pU�	YE��b_�ª�B�#qF`�WRp��_�YD������VFRIEN�D���UFRAM�δ��TOOLȆM�YH����LENG�TH_VTE��Ix���[�$SE�`~��UFINV_�@��5aRGI��N�ITI���XX�l	�J�G2J�G1T� U�D�d�u���_Â#O_p�py�ၻ��"n�C	�zŔ�C ���ʖ �G��zr2�� @ 9�qC����d�wu��ysF� ����p��X n#�E_M�pCT^��H��f��<u6�	�G�#WV�z�G���Dh LOCK~�U� �������$� �2���~�D ��1T���2��2�3��3���:����V��VP=�"�=�F�V��!Р��/������p� xṿ����Prƻ���������E����؅�!��AC�PRs�!�}�S���`���r
��a� 0 5�ؠ�V��ؠA���	������
MŽS��� ح�R��qda��$RUNMN�`AX2q��A���L�+"��THIC�x� w �u��FEgRENg���IF���x���I����V��G�1&�*Ԅ�1ٲ[�nI�_JFR�PR���
��RV_DATA�q� RD�[- 
�AL� �x�Α �b{�  ?2� �S��`?�	� �$ Z="GROU��!�TOT����DSP>��JOGLIYs�'E_P�PrO��\�7`��bvK�p_MI�R�.䎐MQ�O�A	Pp��E<�o��t���SYSE�ib��PG���BRK���v$ A;XIa  �⃃����Ҽ�A����H�B'SOC��T�N���{16�$SV1��DE_OPNsSFSPD_OVR4 ʓ���D� �OR$+��PN�P,�F��,�6�OV�SFa���d�$�F}�ja2㒓���ҁibLCHH\R�ECOV�n��WbE�M����RONs����_���� @��9�VER��n�O�FS9�C�Я�WD�E���A����Rh��T�RBq6aY�E_F�DOh�MB_CM4kS B��BL��.�u��8�V摁��p�d��]�Gv��AM��`i ������_M� �[r�ec T$CA���D��HB�K�q�vIO��8,�a��PPA L�1\D��bDVC_DB<���q�b���ja�1���y3���ATIOi`jqcp�U�� �efCAB�����J��������__p�vS�UBCPU�b�S v��`_��p"�`'}����b"�$HW_AC� Ip���'ɣAx�~���$UNIT���� � ATTRIx���"�CYCL���NECA�Y�FLTR_2_FI#�0�h��f��LP$����_SCT��F_Ʋ'F_�,E2�*FS8�a��"CHA��-7p�1�Pr�2RSD  `�b�����a�`_T��PRO�MFpEM�	`_���Ts2��c s2���5DI&�~�tRAILAC���M��LO�����5��������P�R�S̑{�dAC�p	��FUNC!��RIN됫�|��@�DEqRA�@�� ��C7`�CWARB�	BLƑ�G�DaA�K�!�H�HDA��0�AX�C�ELD�p𐒡@S���A�@STaI��`U�ѓ�$<�gRIA�q�bAFQ P=��S��U �����3MOI� PD�F_ꀔ��qHpLM��FAE�HRDY.]�ORGEPH�0���|� P�UMULSEP���`'���0J(��JC�X�S�FAN_�ALMLVBs_aW{RNfeHARD����v�䐟p�@2$SHADOW��0��a@�b��_`+q�ї�_���vAU�Rx4\rTO_SBR��e����j� ��A	sMPINF���!t6Q'sgREG���aDGBPb��V�p.�l�FL�%!���DAՀ_��P�CM��N�YƧB �V  ��� �]���$N�$�Z�� �Ҭ����7� �|�EG���ӌ��qAR��#��2p?��wP��AXE��wROB��RED���WD���_F���SYм�!���h�Sr�WRqIE��v� STR��(�`��7�E�!�����a��B����@C]D� OTO7q����ARY����.A�̟�#�FI��9�$�LINK�Q���Ry�_���6��N8�XYZ�bB�7P�'OFF
 �7�+�%�B��yB�����0}@��FI� ����h��yB
�_Jဓ�5�����`Ȅҋ8���H�TB�b�CL0x�DU �9AETURa`XgSW���brX���FLz�@��#�pu�Y���3\���� 1��K�M����31�DB`%8��`'2ORQ�6�� �C��}�DB��>��P���%�����\q:�OVEA���M90=ѻs[��s [��rZ��`X��aY��  X�O�~@91�P��B�F� ���=�S�B�_���s�����ER�A	BEBE��� QC"�Aб�����E�2��Q&QAX���Q� �! �|�A��+a����� @@��O���n������N���1����`��` ��`��`��`��` ��`��`��`�!���� �Rg�DEBU�#$�A�c�2���3�ABGE�;�V�" 
�Ҷ�� �z!$�
�$��$�@A $�O�$�n�$��$�N���T#��R����LAB⬒�� �GROh0��l� B_�1 	ƞ�>��`����8���a	�ANDàE @��<���aF� ���q��Z�Qi�� ;�NTq`�cR�C�1=���
�� �pERsVE���p� $q�ڱ@A�a!��PO �`X �����Q�p��p$��TREQm�
��Q����ƑR2�oP@_ �� l=���fESRRҒ�IV�����gTOQ����L�%��Ď�z�0G��%�%�"��?�!P � ,��2 뺱R�A� 2� d��D�p�  ��p$O��2�Pvµ�OCQ� �  }YCOUNT����FZN_CFG���� 4� ^v2T��d�"���m W k!�E�s� ��M �08b�����X��0�CFA~P���V�XA�@�����0���O rA�P�b�pHELkp~N� 5ސ�B_BAS�#RS)R]vm@;�S�!YQRB 1�B 2e*3e*U4e*5e*6e*7e*98�5!ROOGP� ��:�NL�q)�AB���@C ACK�I%NT80�sU�``x1�)_PUA��b�2OU��P�@^x"#��y0��b�TPFWD�_KARlfpZR�E���PP�&Q�@QUE]zROB�2����`�aIb`�"#8�$C80Bv8�SEMա�6t�`A�STY43SO�0�dDI1�@pr�1aǿQ_TM�s�MANRQAF8�E�ND�d$KEY?SWITCHS3h1�#A�4HE2�BEA�TM�cPE�pLEPks1���HUg3F�4�h2S(DDO_HOeM�PO�a� EF"�PR���rS����v�@�OaX �OV_Mx���`pPIOCM$���7��##HK��q� D5�_w�U��b�2M�p�44�%�FwORCcsWAR�R�9WOM�p �� @��˓�`U��P��1�V2�V3�V4���Ox0L�R�<�^xUNLO.0�d�dED�a  ��$$CLASS� `���.a-�&-� #`S�0+hw9`��?a�IRT?�,o>`AA{VM��K 2 je� ?0  �55a�o2�h�o�m ��jA	�m-�k`��o2v7u�lV}b�a`h���t{`BS4�� 1Li� <��� � 2�D�V�h�z������� ԏ���
��.�@� R�d�v���������П �����*�<�N�`� r���������̯ޯ� ��&�8�J�\�n��� ������ȿڿ�����rC`�AX�� `û��s  �%�I�N.�@�$�PR�0X�EQ�}�`�_UP$MIl�ja{`L�PR� ji`��tLMDG6P�g�`��P�IF �k`d ��0�B�T�b�߅��ߩ߻���, 
 ���n��o�0�B�T�g�x�������yNGTOL  �{�pA   ��
�{`�Pd�O ��� ��=�O�a�s�6b � ��u���2b������ ������&J4Z��������� �*<N`r���zPPLICAΗ1 ?je}�����Hand�lingTool� � 
V8.?30P/58��
88340���F0!�755�����7DC�3�����ޝ��FRA� w6*-  !�� TIVqŵ>�2�#UPn1 ��\�}PAPGAPONf`��.za� OUPLE�D 1�i� �/03?E?W?�_CU�REQ 1�k 	 P�a7a<�P�l�?p�d}��33b9b� ���4H��522�:HTTHKY�?Kx�?�?ZO�? 6OHOfOlO~O�O�O�O �O�O�O�OV_ _2_D_ b_h_z_�_�_�_�_�_ �_�_Roo.o@o^odo vo�o�o�o�o�o�o�o N*<Z`r� ������J�� &�8�V�\�n������� ��ȏڏ�F��"�4� R�X�j�|�������ğ ֟�B���0�N�T� f�x���������ү� >���,�J�P�b�t� ��������ο�:�� �(�F�L�^�pςϔ� �ϸ�����6� ��$� B�H�Z�l�~ߐߢ��6�s5TO��/�#DO?_CLEAN�/�$�6�NM  �� a?��������g>DSPDRYRL=�p5HI� `�@q� 8�J�\�n������������������m8MA�X�����17.X��-!*2-!�"PLU�GG0�*3�%PRUC��B^�b�'���O���
�SEGF� K���^� p�8J\n���LAP�(�3�� �
//./@/R/d/v/��/�/�/�#TOTA�LPy	�#USENU"; �8?�2�s0RGDISPM+MC� o1C�@�@@
�"4O�5� 3_STRIN�G 1	�+
��M� S�*
~�1_ITEM1�6  n�-�?�?�?�? �?OO'O9OKO]OoO �O�O�O�O�O�O�O�O�I/O SI�GNAL�5T�ryout Mo{de�5Inp?P�Simulate�d�1OutQ\�OVERR� �= 100�2I?n cyclEU�1�Prog Ab�or[S�1;TSt�atus�3	Heartbeat�7�MH Faul<�W�SAler�Y_  oo$o6oHoZolo~o�o�o �;� �?�o�o);M _q����������%�7��oWOR� �;o��oI����� ��͏ߏ���'�9� K�]�o���������ɟ۟�PO�;�Q� ����6�H�Z�l�~��� ����Ưد���� ��2�D�V�h�z����DEV���*���޿� ��&�8�J�\�nπ� �Ϥ϶����������|"�4�PALT�m [ч�5߃ߕߧ߹��� ������%�7�I�[�m�������I�GRI3 �;��s���'� 9�K�]�o��������� ��������#5GYk��� R�m�� }���%7 I[m��������/�PREG_�H �!/o/�/�/ �/�/�/�/�/�/?#? 5?G?Y?k?}?�?�?�?~]�$ARG_o��D ?	�����1� � 	$V	[
H]
G�W+I�0�SBN_CONF�IG 
�;IQ�HRCACII_S�AVE  T�hA_B�0TCELL�SETUP ��:%  OME_�IO]\%MO�V_H�@�O�ORE�P�_�:UTOB�ACK�ASM�FRA:\5+c _5&�@'`�P�5'dX� q^ ,H5-�_�_�_p�_�_*o]T���0o Xojo|o�o�o�o5%Eo �o�o&8�o\ n�����S� ��"�4�F��j�|��������ď֏�� � PQ_3S_\AT�BCKCTL.T�MP XLED.GIF _$�6�H�Z��ZqsAkA0P�INI^��U[E~-SMESSAGw@����A�0��ODE_!D�@zFDV��O��ǟ�-SPAUS'� !���; ((O �2�1��Q�?�u�c� ���������������;�I����TSK�  
�d__0PUgPDT����d���ԖXWZD_ENqB��WJ��STA����1���1WSM_C5FO@�5]E�7~�GRP 2�� 	BB�  A܊��9XISI@UN�T 2j��C � 	z���A���Ϭ� ����	���-��=�c�nf�MET� 2u��PNߧ�J���^�SC[RD�1��P	�EB��$�6�H� Z�l�~�]_5*Q{I� ��������(���L� ��p�����������1�k��73QGRn���蟬	��NA�@�;	�3T_ED��1��
 �%-��EDT-���J�L�U /dD�@-3Sz5*,B&o�Fs^&  ��2 �K�wʹ�E��	�-3�X5/ |�/|/��k/�4�/$/?H/��/@H?�/�/7?�/5�? �/�??��?O[?m?O�?6LO�?�O�? �uO�O'O9O�O]O7_�Oe_�O�A_�_ �O_�_)_8�_�1o��oxo�_�_go�_9�o o�oDo��oD�o�o3�oCRS_���] ��Ug��	 V ?NO_DEL'�GE_UNUSE�%IGALLO�W 19	��(�*SYSTE�M*��	$SE�RV*¯�Ȁ�RE�Gх$��ȀN�UM���	�PM�Ut���LAY��Я�PMP�AL��J�CYC1�0U�h�R�V���ULSUH�
�j��Ӄ�L��ݔBOXO{RI��CUR_ʐ~	�PMCNVD��ʐ10~�0�T4DLIȰß�ˋ�$MRߎ�&� &�ϲ����̯ޯ����y	 LAL_OU�T k��(W?D_ABORo����m�ITR_RT�N�����m�NONgSTOM �� Ը�CE_RIA_IT������˰F�ѣU�c���_�LIM߂2`? �  N��NϢ��<��m�`����� ?Ϡϲ��ϯ�
�����p��PARA�MGP 1U��Ύ�O�a�s�2ܟC>  CV���f���z�ߵߗЇ�Б��Ж�Р�Ъ�д��Ԛ٢���������C}���ǀ Cїе�+���?�ɲH=EC�ONFI�w�nE�G_P�1U� 49��������������E�KP7AUS�19� ,�uG�Y�C�}� g��������������� 1U?e�!��M��NFO 1v(�� �=����� �	̀���@������%^���A�f��� D���D�q}D�Q�6��p���h ˰O����ǩ�COLLEC+T_�(��p�EN`���\�IN[DEx(����!�1234567890����H����H,��)'/ L/�|&/8/�/�{j/|/ �/�/�/�/?�/�/? e?0?B?T?�?x?�?�? �?�?�?�?=OOO,O �OPObOtO�O�O�" � ɶI�O "������O_a_s_�_WTR��2#](�8Y
�O�^P�$,]�Z��^Y_MOR"�%� �9�Fe�Fi^oLo��opo�o�kb�#�&-mB�?>�>����aR�Kt�A�PMy(���a�-=� Oas�ϗ������^@
�����` *c�PD�BO*���Ecpmidbg�C����U�:��ii)�p�/���S�  ����e�-�̏���ܧ�m��v�������9��g�^�)�	��fM���w��>�@ud1:˟����Z�DEF )�o7S)ߑc�b?uf.txt��M�� �p_L64FIX +�Q��� ˓�د��ɯ��2� D�#�h�z�Y������� Կ�ſ
��.�f�x�__E ,� ̀l�~ϐϢϴ���p�I�M�C-�]��6���>���=L�͖��MC&c.�Sd(F�'�%d/5ݤ`t��v��B!!������@�߹���>�T��g1�\�D�y**�~***�}��`U�kx*��CÇ�鯇�BDw�4  �E	�a�Ee�3�Ec��Et� �F�3E�Ś�F�B��F����F�YfF�%� G�� G	�߳H�3�y?��  >�33 ;s���a�v  nf�:�q@�a5����b��pA�a�t�<#��eDQ��7���F�RS�MOFST 'X�f�G�T1#`DZ�-2!���
�*�;�0�R�L�?����<�M��T�EST�0��FR�z3SMx�C�A%�z�*e����| C��B��C��pn���*:d��b2Iy4<�2T_�PROG ,k%^�/%P�NUSER  �1��KEY_?TBL  -e1�]�(��	
��� !"#$%&�'()*+,-.�/�:;<=>?�@ABC�GHI�JKLMNOPQ�RSTUVWXY�Z[\]^_`a�bcdefghi�jklmnopq�rstuvwxy�z{|}~�������������������������������������������������������������������������������͓���������������������������������耇�������������������s���A� LCK#xD#STATi/�0_AUTO_D�OG㺒�+INDTo_ENB�/ �"���/�&T2�/6S�TOP�/�"SXC�� 25K�p8�
SONY XCg-56Q{��p_�@��͞b �P�АX5HRC50�z-tx?�>7�?�5Aff�:�O"O �?GOYO4O}O�O jO�O�O�O�O�O�O_�1__U_g_�\TRL�� LETE6 ��)T_SCREE�N -jk�cs��PU0MM�ENU 16� <O\�o�u�_ oIo��&oLo�o\ono �o�o�o�o�o�o 9 "oFX�|� ����#���Y� 0�B�h���x���׏�� �������U�,�>� ��b�t�������П	� ���?��(�u�L�^� ���������ʯܯ)�  ��8�q�H�Z���~� ��ݿ��ƿ�%���� [�2�Dϑ�h�zϠ��������b��S_MA�NUAL"?�QDB;CO� RIG�Ws)�DBG_ERRL&� 7�[���������� O�NUMSLI I���dD�
O�PXWORK 18���&�8��J�\�n�DBTB�_�Q 9<�����K,�DB_�AWAYW���G�CP D=����_CAL �/��S�Y!0�UD H�_q� 1:
����0,R0�T�P�A�~���_M� IS� ��@� ��ONT�IM�W�D����
2#�MOT�NEND'"�RECORD 1@�� �����G�O�N<����z�� �G��Nr' 9K����� �����#/�G/ �k/}/�/�//�/4/ �/X/??1?C?�/g? �/�?�/�?�?�?�?T? 	Ox?O�?QOcOuO�O �?�OO�O>O�O__�)_�OM_8_F_�_�N�ex�_�_�_<_�_�_8�_'o�N�U(o_o�qo�_�o�o�o�o�NH�I�o�o9$82o�N���p���(�����N���_�K�]����TOLERENC��sB����L��O��CSS_CNST�CY 2A~� 	h���Џޏ��� �&�8�J�`�n����� ����ȟڟ����"����DEVICE ;2B~� ��r� ��������ϯ�����)�����HNDG�D C~�Cz�<���LS 2D\�;�����Ͽ�����=���PARAM E/���?�)����SLAVE �F~�J�_CFG� G/�)�d�MC:\��L%0?4d.CSV(��c����A ��C	H��n�n�)��=�
[��)�-�Z�j�X�<W��JPъ�C��_CRC_OUT H��<�+ϑ�?SGN I�����\�17�-MAR-25 �14:49��)�05��6:01����� Ze��7-�)�)�*���o���Im��P�u�G�=��VERS�ION ���V3.5.20���EFLOGIC� 1J% 	���* ������PROG_ENB�����ULS�� �,P��_ACCL{IM�������7�WRSTJN`����)��MO��
��x�INIT cK%
��) v�wOPTp� ?	�����
 	R5�75)���74��6J��7��5��1�2���6����TO�  ��@���V.��DEXd�d��x���PATH ����A\����IAG_GRPw 2PI�|O��	 E7� E�?h D�� C�� C ��B���C��n�k�����C���Cm�B�N��BzoOB�)��Bk��f383 6789012345����B�  A���A���A��A�O�A���A{+A�s�Aj�RAbJAY%, x�@���p��G!���A�����BA4h���x�
"�����"�Q�A����A���A߈��A�� ���hAx~�Ao��7Af9X��?$>��mF/X/��h�����("_�AY��;AS�TAM��^AGdZA@��A:bA3�%A+�-A$���)�/�/��?�*�@�;d�6����@{�@u�-�@o�@i�7�@cC�@\�j�@V{N?\0�5�?b?t?�??@_���@Z^5@T���@O�@IG��@C33@<��@6�+@/<@(�`J?\?�?�?O��8s� nE�@h��@b�!@\��0Vff@Pt@I�hs@B��@;�bOtO�O�O�O�' 6]^_p_N_�_�_0_z_ �_�_�_�_$o�_�_
o lo~o\o�o�o>o�o�� C"�!30�2KA�@^�>8Q�r��R�?�  *u^7��ŬFr'Ŭ5A�FRu^@�p��nv�@@�pppE�@�[ Ah���uC=�+<��
=T���=�O�=��=�<����<�p�q�xG�� �?� �C��  <(�US�� 4jr�D@���Y�"�A@w�?f �oX��mf�������� ��ԏn��
��.�@���i?#�
b���\>�pn�^��G���G�^x���R����^8�ۑ�5����CnB��L]_u��&�
P;�'f�d��aQ�{���dD�  D�  C΍��̯ޯ 8����@V�ǯD�ïh������3+��Q�ҿ���� ��,��P�;�%ZN��Dϥ�CT_CONFIG Q-y��#�c�p��� STBF_TTSd�
����C�tV����MAU^�����MSW_CF���R-  ]z��O�CVIEW�SY�i�����߽��� �����G��.�@�R� d�v��������� �����*�<�N�`�r� ����%��������� ��8J\n�� !�����" �FXj|��/�����//j�R%CR�T�e&�!�,. V/�/z/�/�/�/�/�/��SBL_FAULT UI*n�1GPMSK��$7���TDIAG V���e�2�UD�1: 6789012345�2��?�P�Ͻ?�?�?�?OO )O;OMO_OqO�O�O�Op�O�O�O(� �>��;�
�?%_��TRECPZ?l:
z4l_?� �?�_�_�_�_�_�_o o0oBoTofoxo�o�o��o�o�o�O_/_U�MP_OPTIO1N��>*qTRR���:!9KuPME��>�Y_TEMP  È�3B���p�A�p�tUNI�7��şqF�YN_B�RK WY�)8E�MGDI_STA`�u&��q ��pNC�s;1XY� ��o7�*�~y���d ���� ��Ǐُ����!�3� E�W�i�{�������ß ՟����r�,�>�P� b����f�������¯ ԯ���
��.�@�R� d�v���������п� �����%�7�I�[�u� ϑϣϵ��������� �!�3�E�W�i�{ߍ� �߱����������� /�A�S�m�w���� ����������+�=� O�a�s����������� �������'9Ke� [������� �#5GYk} ������ /1/C/�oy/�/�/ �/�/�/�/�/	??-? ??Q?c?u?�?�?�?�? �?�?�/O)O;OMO g/qO�O�O�O�O�O�O �O__%_7_I_[_m_ _�_�_�_�_�_�_O o!o3oEo_Oio{o�o �o�o�o�o�o�o /ASew��� ����_��+�=� WoI�s���������͏ ߏ���'�9�K�]� o���������ɟ۟� ��#�5�O�a�k�}� ������ůׯ���� �1�C�U�g�y����� ����ӿ���	��-� ?�Y�c�uχϙϫϽ� ��������)�;�M� _�q߃ߕߧ߹���E� ����%�7�Q�[�m� ������������ �!�3�E�W�i�{��� ������������ /I�Sew��� ����+= Oas����� ���//'/A7/]/ o/�/�/�/�/�/�/�/ �/?#?5?G?Y?k?}? �?�?�?�?���?O O�?K/UOgOyO�O�O �O�O�O�O�O	__-_ ?_Q_c_u_�_�_�_�_ �?�?�_oo)oCOMo _oqo�o�o�o�o�o�o �o%7I[m �����_�� �!�;oE�W�i�{��� ����ÏՏ����� /�A�S�e�w������� ��������3�%� O�a�s���������ͯ ߯���'�9�K�]� o���������џÿ� ���+�=�G�Y�k�}� �ϡϳ���������� �1�C�U�g�yߋߝ� ��ɿۿ����	��5� ?�Q�c�u����� ��������)�;�M� _�q�������!����� ��-�7I[m ������� !3EWi{� �������/% //A/S/e/w/�/�/�/ �/�/�/�/??+?=? O?a?s?�?�?�?��? �?�?O/O9OKO]O oO�O�O�O�O�O�O�O �O_#_5_G_Y_k_}_ �_�_�?�?�_�_�_�_ 'O1oCoUogoyo�o�o �o�o�o�o�o	- ?Qcu���_�_ ����o)�;�M� _�q���������ˏݏ ���%�7�I�[�m� ������ǟٟ��� �!�3�E�W�i�{��� ����ïկ����� /�A�S�e�w������� ��ѿ�����+�=� O�a�sυϗϩϻ��� ������'�9�K�]� o߁ߓ߭��������� ��#�5�G�Y�k�}� ������������� �1�C�U�g�y����� �����������- ?Qcu���� ���);M _q�������� �	/%/7/I/[/m/ /�/�/�/�/�/�/�/ ?!?3?E?W?i?{?�? ��?�?�?�?/OO /OAOSOeOwO�O�O�O �O�O�O�O__+_=_ O_a_s_�_�?�_�_�_ �_�?�_o'o9oKo]o oo�o�o�o�o�o�o�o �o#5GYk}��_ �$ENETMODE 1Y�U��  �P�P�U��{��pRROR_PR_OG %�z%�V��&��uTABLE  �{oe�w�������rSEV_N�UM �r  ���q���q_A�UTO_ENB � �u�s�t_NON΁ Z�{�q��_  *����%����Ā+�*�8<�N��HIS���Q��p�_ALM 1][�{ ��T��P+O�˟ݟ����%�S�_����  ��{��rj��pT�CP_VER �!�z!�5�$EX�TLOG_REQ�k��ቼ�SIZ\ů��STK�������TOL  ��QDzs��A= ��_BWDJ���؆K�ԧ_DI9� \�U��t�Q<�rU�STEPa�s�|�p��OP_DO���qFACTORY�_TUNk�d̹D�R_GRP 1]�yށd 	e�#��p��x����� �n��So �k� ���W��i� z�dϝψ��Ϭ����π	����?�*�c�N�@�� @畱?���@Q�j�?
 E���R���j��xd����E7�� E?p D�����L�D�%��  �C���K�B�  >;�  A@E�o�o@UUUc�UUo��&�>�]�>П���ި�E�F@� F�5U��{�L����M��J�k�K�v�H�,�Hk�{��?���Q�9tQv�+�8���6h��%7�{�W> �O���sO���Gj ,k���rP,�FEATU�RE ^�UK���qHand�lingTool� �� rodu�Chinese� Diction�ary��LOAD4D St���ard��  ND�IFAnal�og I/O�� � d - ��gle Shift���F OR��uto� Softwar�e Update�   J70 m�atic Bacwkup��art �Hground �Edit���70�8\��ameraz��F��D pr��nrRndImMޤ�PCVL��om�mon cali�b UI q.�pc�nf� Mo�nitor��ws�et�tr��ReOliab	 ��jp �Data Acquis������ Diagnos�D����� Doc�ument Vi�ewe���
P�C ual Ch�eck Safe�ty� act.�Enhanc�ed UsGFr�w ��\weqpxt. DIO � �fi+ t\j7�endxErr� L*  � �{'s  ��r��� :���T "� F�CTN Menur`v���t I��TP In�fa}c%  48\� �G_ p Mask/ Exctg�� �o��T Proxoy SvH  5�p��igh-Sp�exSki� "� #1��#�mm�unicC onsn�apd�!ur ������"con�nect 2Pd�in� ncr sgtru�� I �KAREL Cmod. LE uaG"�t\ia�%Runw-Ti�Env�z�"K�el +G �sE S/W�?Licen��[�GER  �Bo�ok(Syste�m)�� R5� M�ACROs,x"/gOff� �Pa� �MH�- �: \ac�1MR� �)���MechStop�V!t�  ��0i8���Mixx��dE ��
� �0od
 �witch��Lo�a� �4.�6 k� G�1�3OptmpUHM GGW filG҅ HF��g�' p�mfO Multic-T= i�4pa�PCM fun�'�{3M"Po[�D zQV�HRegit0}r�   mpo� �Pri@F�K _�fcs W g Num Sel�5��� |DS� Adju� P���`W
 4 S|XtatuQ/bUC��� RDM �Robot��sc�ove�� cctNO Rem�0�n��<�SServH10@�#CTXPSN�PX b<2�� "�K9$`Libr����564@e�� X�4H`ZUSoY0t �ssag�E�~� �"�1�VVLO�b/}I- pc
�`�MILIB�mchy1o Firm+p�8� �b"Acc` <hXcTPTX�;��<� s Teln�0�m�}B��5��4Tor�qu
 imula��}�Tou7@P)a51��m�T_ ��QC&V ev. o�cleUSBg poU � iP��a@WdUSR E�VxP+Unexceptx�P�D{D,{f}VC�r�"�"�2�sVD��j�cV��Hk uifoV�S?P CSUI�k���XC�6X`We�b Pl�V��9pjxăa�+64.f���^ r>�T�v�
J�57À�vGrid��Qplay 76� (��`L&iR�;�.��K�\0ARyC; 4 120i��>L#AsciiV!eRpDAG�d��UplE@x��� �@CollW�;Gu�� of^QޝPI   1�s� ���t�0t8FK���Cyr�p  2*Porie�  ld�aFRL��1am͉ RIN�T��MI DevfO0 (&ax2 ,�0<�%(}t\rb�A/~��Passwo���:O" 64MB� DRAM�

!� 0ڢFRO�q�G`��rciPvis��y6BW�Wel�ds cial�4 )��ell���!P�shK���wmrEwd�cXE|�( p�v�� wmd�ty	 s�PRa��P0�t!1m@.
)�8�D�P����X�P+�D� 2b a��@�r�dr�Pb� q�D�rT1� egedv� OL��Sup�rx�AR8sOPT "W� ! � d��; cro�V  �SHe�[�  ��
gq�<�u�est;`LO SS���e�tex 	E�$`p$![b�Us�CPP@ �4YPVGirtW�St�e~��Pdpn�x��  �� SWI�MEST f� F�0���ui.� &���ߖ� аߞ��51 J����(sFr�ߕ�II)����on��!���M!=���	QY���f>�t���mfV��լ���Ҍr ���?���&P�3����Ҭb9���eie�߽�n\p���\R���ҭ`A��2�p�����!
!����O<����7 J5�����5�ӝ1Q��\a�r7���XPR���k "��}��b���r�`P���lnko�0���`1��RMJ�Ո��;���M�����Hs54���j883�]DER�N��Ffh�M/el���չ1d/������d0�/ ��|B�/�( �/��<���/��p����.fd��/��ASTC?��6�16�/��g HS0|?z��as���� ��1��?��0�?c�r W$O��!`��%�rzP]O��t\aw xOV4�`�O�$�a�O�Ҁ���O����O��.E�N _�D�`<_��itye_?��v t_f�� aO��IF{?p�Ԉ`���) "s_F�Epa�O-�>n1!ONt.vTo5!�_���F���o^837�o*QogW-���o�/p��X@�PDT4���_��ze�OHf4L�_\79���MN�`�����f�tro�9?6�x�i0���J5!9L��%����Ak��P����_p�o�Fp�_-o�@�?(�f91'?�pm_d��O���ٟ�O.�pe����m\�A��/_8����2.p�͆cW_�֮͠c�a/�\ R8���(Las$���O_���0x���bo��<����I�̿"% ���K��/?�sif<Ϟd�?�3NT+���Se�� ��//�C/�����'337��iUf\�����$SG��Ԁ6h��RDYLS߱�oI��omw��_#�ps0 �����hVmj��93����E�ogW�P��ch\?�I���ퟓ� �o����rv	i7�]S�/������V(st,��F���&@�tl�u&5/�$���T
�hWi��ݶ�Se��6O��sr���	��! ��y8P`�dr׏�o3'PRI���a�O��/	X/��spr0�ߕ����Li?/���3 H6x/�d94�'��63�q54 H��/v653�/r4 	H���&0�/�'��� X?v72�Ie?&�g13;?��7�/5�8r?�'6�/��Lo�_��t �ͅA���Oc�m�osK�!����O����,�O9��O�ONS�ualP_��8�?�a_?�8�_��w9r+��j83�?!��_]���NDSO-�fd7O=�!�Y�ad�O�9kl�o�s_#1 �o��ip#�-Et�op�gRIN,��/I��f��VA�=SE_���0
S���Zs 0+ͅcmg��Z�� 4@�"�ut@[/�of��`�M�r�p���@����596O_��4Џ��U��#o(�1 I�c5%r_����e`���G�������8c��AL"����lg33_U�oy� -<�t
��	e�@t���RTU���h�0z�xo��vo;��'O�52 ����4���'�Yu\�� vOAȳ��4I`FĿ
d -d�ݕE��� (o��[�"E3�yo��W�el_��������WMG�Ϣ3aP@�Ϣ3wmg[����߂�c- ���On�45�?��fCMk�IO��  �ߪ������1���2�g�y� R�;�3Co���4(S�`�`⯔�Ġ��3IF����� !(�z�0at���NT��q���Ra8��i5᯳W2\��� O��W?��˿�ݿ￘��7��4Si�Z/<��=�K�!�cl��i5\sw/�S�A�D���CVt�Dt.�Q�mt�_�e���V�-V�  /6��N#lo��1��\�O�/C �/�4 �/��i�e/�/1_�W62d˟��o�/�eJ7���erv�?�) 9"�?�svh�?
o0�N� �?�.p[�t�vhmoO�U749�LOR`r��OutIlO?�t\�?��j�_��//�/h_ mp�c��y�9\KO�j`�_�/�_�uXP�/�D�H8gO}�oOnn�O�%N�߬u�'o���n]`���oRCM�o�un�_��$./�_#��m  H552��abe�q38BS�R78�p�q�r0���libJ6�14�cATU�P�@rmc�p54]5zPsgt�r6��VCAM�3�CRI�p\rc�pCUIF�  �q�2�ptd.f�N�REN rco�p6�31  - Pr�pSCHV� Di�DOCV>aI]FL�CSUJ18��0�p1}�EI�OC  ��4�p5�4�pR�`4�9�pg�m�SETf�Sta��q�qlay,�p7��q�0MAS�K�SPRXYVZaap�7f�C�pOHOCOC��3.3l�r�p\c΂51�p���qapp.�q3�9f�j50�q�u;st3�LCH��A`
OPLG�1�"�E�� "L3�M�HCR  08 u(ĀS@�Reg��CS�p�1H��p��q�5�p08\�pMDSW  URGw��MD���sOP��\.!�MPR�ra�4��Հ!�o�f��p! p���PCM�H��R=0БPath���p�@aH�ՀRm����pT�P���Հ816�5�0�pg��āS��o�l,�9Ղ:�FRqD�p(Q�pMCN���cc�H93�pL{NP��SNBA@��rSHLB��֑S�Mx�lrn?�63��p��q2�pL�HTyC�pX�TMILVs0�r�T��PAu�Y�msȡTX>aEN��[ELU�th��0�@`�8�qHѰr9��`�ρ95�p �Հ7UEV��adi�n(�C�����pUF�RI�eeO�VCC��pt�VCOY���V;IP��spd�[�iI^�p�X͡tsπ�WEB�p��?�HT�T�p L2�R62n�pCoo?�CG���d�IGt�
P�RI��PGSN n�g�IRC��ne� ��H84�prd&6�R7��@�R��L�{53�p\lcl�q�8�pD" #4�6�M� ��52�8�R�659��|�5�r� dK�6��p��4�4�9�YpS��p5�̰L�0=6�pVG MD�o�7g, ��66�p���ðAWS�pJ643�LIက�V��pczdҡ��u�GD�����q�%�h�TY�� ����TO�p<q�q6��g��|� �-@��OsRSY��R68�p�3��OLp�ģOP�IɰsguK�SE#ND�/аpLP�T�qS��y��ETSɰ2!�6�U����-�o43 !D�VRu��ry:�IPN��o�nF�Gene��o{aytD (S��E���I�0�֙���p��ytt\sg��g ="�ր6h��L�yt\str�ոA��<�A��hk_t���yt����es�լr��{j7��mon.��(�A��d@6��s-@����yt46\�`Q����qh3��zDlli�4�F�lc�`�$rt{���¥���yt��w�x�U�Ӑh8��nde��AxV絰�����N��ͰH��epCen���yt�T�ՌĢ��ob3攢��hS89����p��Pv�sed����4 J7/R805��0l���:�`"t644������ II���r�p����"S��/л%���594G�tomt���!�R J�ؖ� ��Se3�ar3�E�t32�%�QsysG�F ���������etr��ur1nk����20�xc78���'�rn6������\jtET��
jo��ta.C����gr������`� ���<���ge�.��017��2�ytL�yt75b���Lj(t���7 "P��T`dc��) ���	����r��1%a�t�@O���p��daW(?�4tv/ 4oh��c8}���s?yR�?��=logm�?�;ild�?1<d�?N�@ ���0@O�M���p1|O�;x@���ytV�B�1���O_�	8�7aicC 2�9���C��7��6o�E �� `�E?kedg?y=wm�`ORhl$_�2G&�he>�m_��7�5�l�O 24O Oaw�4OJmdh\o�;dhq2���osqz�o�kl���o�o��:��+�F�et�'-�6J�8"WQ��1 (F����pDa�0��f�r{F� �� �f22�.f�FusS�pkYg�M!INgD�x���,��u��o�{Ώ�522�xsiR=C�n VM��^��992�W� ��J9�b�st�'T��Oo 92\�6CMR/@d#Z��O;��ݎv'�D��tmF����f8��vat��t+9�>e��6ft"/��zC_v(��ɟ?�4o ��,���կK����cvsw�8��Dni�o��lb��蟮������W�\���vsmTڴaz�"����ο��of���1ow�(ώ�slw���f���e�w�����*ԣvr�ys�+N3Ge�N���Y25:�oa]d��(Na�NJ�?��nd�� "N�wV  �(F89���rrd�6`��le&���C�U�14;��Ok7\��8�b��rk&,��gl���P��g�Gt��il�������  � P2^���38��r �����0��J614~�ATUPj�N��545����6F��VCAM��/CRI!7� , �UIFB���2��a{ns��CNRE�'n��631��RI���SCH�u65oDOCVN�ns� GCSU�T|���0��~HAEIOC%� "��54��R6�965\� ES�ET�W�����7� Cu� MAS�K�t 1P�RXYUJ N 7ܺל�OCO�om.�513r�,,���x��� ��98\t��X��]�[39�v!����oftwL�CH!g�OPL�G:�950aip�P]P��e f,eS�r��CS��x���g_lo���5� �pDSW�6�r70<!Pl �DKOPP4�PRQS01� n A�d����X#PCMAa ��0�%����vdv; �A�
TX��0��1�ADIG� �!�H ,S�r723���9AU�+ FRD�!h#RMCNr	H�93��R2SNB�A"�C+ SHLB��	SMp5�n m��J52�HTC����TMIL6�S�e���PO�0PA��86*TPTX��VR�0ELA4oo�l,��� P��8���\sv���qS7RVT��95Q$�95A\et� U#EV�@a\AC!]��[AFR!r��C�!ol.�VCO���P��VIP�4e��� I�t34[S�X���WEB���@(�1T��,�l�2tQ, G�Eg\-tkIG�E#@`PgPGS"�PRC�4o"TAN��84���#R7�taQR\�(
R53�tR�J68��R66�a52a- E���R65qr I�m�5a��l��5;73R64q�h��q5`M� 061%��BFf�R �  ��WS!40.�ACLIQf9�PnSniKaMS�E��Rn`��597{1T�Y�476 J, T�O��L���6�9 u(k5Pfer@�ORS�CR68���\sn[!L%C;SN� OPI1Tp��\0� ��sn.��L��E �bS�fX�0ETS1T����h#�0�a�P FVR� ��,QN�4�GeneN�a
@�Dx�x���yMG" �y<���yg_cc�y"�xcmg_�y��yGvth�yR�x3(��,�>�P�b��z1��z!� cv�yon T��yh"�xhr�x�b݉1p�`]�iA�y CV�yCP �z��x��xpt���	q�ypse��ܨ���r57� I�n���xy͉576��(p+�)� �����L� "Al��w6\�ab����j8<�B���h ��PR<�J8�zPxC;�8�J��ps��P��x96\{�(P�y�����A�xlY`� -��iv{�oR DM<�H7�z[H6�{66�3�18�x�[�tor��������y�m�!��s�Z�]�2����na�lۺ��)�޸st�K��}str��yp1sk��=�\p����^�xj932|�C��@}�)�x8R�x2}�d����.|�޸_w��.�}hk_k�FH��z�9!�xke*�n�9�5
���yhe�z8�8,�f�l.<��H�et_w�y�"�M�c� �� �zba8k�H�Z�ent��h�\m���s����  ��d�༛�Y�;�(�PZ�@�z9Pf�yv�@ ��.������ l�n��( l�gd��=
iƋ�! Z���+�00iB\�H[�H����� -�h[�C" #���82��2�@}�O�R��� ���iB/�̿N@�"F���f���h@+�=���tk� 3OR����83�i1f�t ˚�~nc+�&�fc����5���835�z����i�;˱5:�B�ri��E�R���b݉ (ˊn�g,�@�,4�*R`ȭY�k�xmo�`�]/��p�+��ptp�z(�5\pk�=O?�A�45[ڈ��0�/�/@ ?S�i�k߽�ij`��
��?�+�db�^�� s50l�a��tx���S�[d G��yϋ�ce��0K�5�0�K1�y�6hu�Je�RDE���yqInt�
 Pa���(�9\g{�H�9�19[�p�\:� V=i��tool<?ވ:	�J[�uppK/=_��vk{��K[��Z� �Z��O�O�O�8�OK�8H��?��_rj;*h��ndr{�H]end$��Ir:�(�3��o�>�73;���/�&7 ;*��{X�j�|����"�4�  am_x�O�ve�ʘ���v$I���o�?|�xj{���� �Tz{�] R�5;�J9�;989@ﭹ���_��p�m
��
�`����e�kR� R�}++R7�J L:;) "���KzR�/p+zx�d	�-��|�	�633�06� S�I~R6�sqt�z��:�LND��7IF K�45��-con{
C9�i�*�ar �jyp�	�d�s "����EN�l�y��s��l�gr括e-����8568��`�zrpi{�x=�H�4 l�^�wnj�! r˛vv�:�nn�}RC:| ��� J9�Z����8[67�13J;6���8 �JT�`��(iR��R|"ٟc  STD���.pLANG(&�����r��ti�����P��q��)0-�� =E��kg
��y`� ��5����R73�0��(��8 (i^��ErrP��,�`���PC��x���rv�ge������8���g�e��a<����	�.ޠ�isio��ck#in�� �R�(���pGi� ������؁��j	��PFK�"��XA��\@��B�P4��!��d��agabbPbbb������P��P��(1��S�P�Р�FS J���J91��685b9!	��02*-4<627���Y��,����X�v��s\�GFSO8����sex��/�vr�����&��v�RG(R68'64����#8	�G (� CCR���I���cc�� �"CkH���9�\�RBT}rgOPTN�4�4�2��4�?�?O"Ocrg�.8EF��8E��
/DPN��d�uD�ion tEnd.qtExa�FINTtER��7tE� ntEa�@�tE�0"tEHQtEhd\m�FHD�F�uD\erh�F���O�A�itE��sF�"Uir�etEhuDtuDrh<�GdCted ����<��n An�U�Y�9p9�Ut2��8��0 E���a�U�`t f�1���2��� m�U�a�U葠U-`s�U�ѠW
 �1����6hޠU R88�U85�1_f4�`�Utia1r�U���it� ��<l"��MR S�f`��fTXP�U��ep�m�f" #1�f!# T�fy��fm�g���e�P�U 2�U 70�Uonjg���@_f� J7�Vipp�fon,�U���X�v4��j79�fc��e]h�98jg�"��\chp�WEN�vd@Pb{'Sto'�� E f�@�VgF0�el�gxѠU��j8svY��f�z��6uharel�UwKARo�Comc�*u�RĆL*wp\ �V�
+vY�u�fp\�e�VAN"���k.�gpcp_f1a!I��[�f4y�wf
! �Gf Co�uar�wf�FІ84_f5� H�fH84�v6�3 H�fH7�v7K79_f24��7rw[69*�65�f1�g�8p��V75�VIC� �f AP7v89�3���R0���B�ecik���Hs�
E8����#fMNS+v�� �VՐ�V�P_f-]�_��Q�VX�\���tch�믅ԠU3\pSfW�T"_fdBe��ZhiYn_� �03jgoX���(ROB�wOG ���AUe�A�^�HR��PxflRuuyQuug�_Sf̉3uh523�.�le*writ�y �6�2�6�5�sv54f�4І40\����H60�v0�h�[�08��+�=��O�a���8< ���6a8v�`��s�75^0��A�rw7��h�����ԕл�3�v3Y�� � �େ20f���� 29#f�p���\ib<f��;s�bs�w��o scbP1oCja��Ly2%�c -k�E"�74�9 wf (W_�	`��3XPF���wvF�E�X�Ϯ`we�Vp�a\wvTf͸�z50+�"WV����֤�u��2�Y �� ��n�te�g�����f04 (�gx��D����'BPXk���I/��`�o�d�@��G��p0v kϥ�ibςhp
om �wfE�A��f��Hfdn���z8�Z�f��ؿ�ra��W�_�oi �<�al��VVAx�V�2�� w996#fVCA��,�vast#/�q� ،�"�dp/fynf:�fi���58��z��D��odif���.e8DP��q (d��o "���o��Rg��d9Ԑ'G��str�S���OAW���wR�73�v16"� R�f�79�2���iT�ra��c�h�/�w�v"TP+v̀��tkpe�c�wor��Z�+RC�59�8��w S5+�809�?��C�f�"z\m�ߦ<����RE���$FL&0�pcuz�6�verv�gsng_��746�_:��S_� Ch�?�� ���8rth��0�897iu3�g���6�f�!��y$�x���� �T����&w& ���rk����`�s�H�VAGǧse�t99�������$FEAT�_ADD ?	�����q�p��	x����� �*�<�N�`�r����� ����̏ޏ����&� 8�J�\�n��������� ȟڟ����"�4�F� X�j�|�������į֯ �����0�B�T�f� x���������ҿ��� ��,�>�P�b�tφ� �Ϫϼ��������� (�:�L�^�p߂ߔߦ� �������� ��$�6� H�Z�l�~������ ������� �2�D�V� h�z������������� ��
.@Rdv ������� *<N`r�� �����//&/ 8/J/\/n/�/�/�/�/ �/�/�/�/?"?4?F?�X?j?|?�?�?�tDE�MO ^�y   x�=�?�? OO%OROIO[O�OO �O�O�O�O�O�O__ !_N_E_W_�_{_�_�_ �_�_�_�_oooJo AoSo�owo�o�o�o�o �o�oF=O |s������ ���B�9�K�x�o� ������ҏɏۏ��� �>�5�G�t�k�}��� ��Οşן����:� 1�C�p�g�y�����ʯ ��ӯ ���	�6�-�?� l�c�u�����ƿ��Ͽ ����2�)�;�h�_� qϋϕ��Ϲ������� �.�%�7�d�[�m߇� �߾ߵ���������*� !�3�`�W�i���� ����������&��/� \�S�e���������� ������"+XO a{������ �'TK]w �������/ /#/P/G/Y/s/}/�/ �/�/�/�/�/??? L?C?U?o?y?�?�?�? �?�?�?O	OOHO?O QOkOuO�O�O�O�O�O �O___D_;_M_g_ q_�_�_�_�_�_�_
o oo@o7oIocomo�o �o�o�o�o�o�o <3E_i��� ������8�/� A�[�e�������ȏ�� я�����4�+�=�W� a�������ğ��͟�� ��0�'�9�S�]��� ��������ɯ����� ,�#�5�O�Y���}��� ����ſ����(�� 1�K�Uς�yϋϸϯ� ��������$��-�G� Q�~�u߇ߴ߽߫��� ���� ��)�C�M�z� q����������� ��%�?�I�v�m�� ������������ !;Eri{�� ����7 Anew���� ��///3/=/j/ a/s/�/�/�/�/�/�/ ???/?9?f?]?o? �?�?�?�?�?�?O�? O+O5ObOYOkO�O�O �O�O�O�O_�O_'_ 1_^_U_g_�_�_�_�_ �_�_ o�_	o#o-oZo Qoco�o�o�o�o�o�o �o�o)VM_ �������� ��%�R�I�[���� ������Ǐ����� !�N�E�W���{����� ��ß������J� A�S���w��������� ������F�=�O� |�s����������߿ ���B�9�K�x�o� �ϮϥϷ�������� �>�5�G�t�k�}ߪ� �߳���������:� 1�C�p�g�y���� ��������	�6�-�?� l�c�u����������� ����2);h_ q������� .%7d[m� �������*/ !/3/`/W/i/�/�/�/ �/�/�/�/�/&??/? \?S?e?�?�?�?�?�? �?�?�?"OO+OXOOO aO�O�O�O�O�O�O�O �O__'_T_K_]_�_ �_�_�_�_�_�_�_o o#oPoGoYo�o}o�o �o�o�o�o�o LCU�y��� ����	��H�?� Q�~�u���������׏ ����D�;�M�z� q���������ӟݟ
� ��@�7�I�v�m�� ������ϯٯ���� <�3�E�r�i�{�����>˽  ¸� ���)�;�M�_�q� �ϕϧϹ�������� �%�7�I�[�m�ߑ� �ߵ����������!� 3�E�W�i�{���� ����������/�A� S�e�w����������� ����+=Oa s������� '9K]o� �������/ #/5/G/Y/k/}/�/�/ �/�/�/�/�/??1? C?U?g?y?�?�?�?�? �?�?�?	OO-O?OQO cOuO�O�O�O�O�O�O �O__)_;_M___q_ �_�_�_�_�_�_�_o o%o7oIo[omoo�o �o�o�o�o�o�o! 3EWi{��� ������/�A� S�e�w���������я �����+�=�O�a� s���������͟ߟ� ��'�9�K�]�o��� ������ɯۯ���� #�5�G�Y�k�}����� ��ſ׿�����1� C�U�g�yϋϝϯ��� ������	��-�?�Q� c�u߇ߙ߽߫����� ����)�;�M�_�q� ������������ �%�7�I�[�m���� ������������! 3EWi{��� ����/A Sew����� ��//+/=/O/a/ s/�/�/�/�/�/�/�/ ??'?9?K?]?o?�?�?�?�?�9  �8�1�?�?	OO-O ?OQOcOuO�O�O�O�O �O�O�O__)_;_M_ __q_�_�_�_�_�_�_ �_oo%o7oIo[omo o�o�o�o�o�o�o�o !3EWi{� �������� /�A�S�e�w������� ��я�����+�=� O�a�s���������͟ ߟ���'�9�K�]� o���������ɯۯ� ���#�5�G�Y�k�}� ������ſ׿���� �1�C�U�g�yϋϝ� ����������	��-� ?�Q�c�u߇ߙ߽߫� ��������)�;�M� _�q��������� ����%�7�I�[�m� ��������������� !3EWi{� ������ /ASew��� ����//+/=/ O/a/s/�/�/�/�/�/ �/�/??'?9?K?]? o?�?�?�?�?�?�?�? �?O#O5OGOYOkO}O �O�O�O�O�O�O�O_ _1_C_U_g_y_�_�_ �_�_�_�_�_	oo-o ?oQocouo�o�o�o�o �o�o�o);M _q������ ���%�7�I�[�m� �������Ǐُ��� �!�3�E�W�i�{��� ����ß՟����� /�A�S�e�w������� ��ѯ�����+�=� O�a�s���������Ϳ ߿���'�9�K�]� oρϓϥϷ������� ���#�5�G�Y�k�}� �ߡ߳���������� �1�C�U�g�y��� ����������	��-� ?�Q�c�u��������� ������);M _q������ �%7I[m ������� /!/3/E/W/i/{/�/ �/�/�/�/�/�/?? /?A?S?e?w?�?�?�?�?�1�0�8�?�? OO1OCOUOgOyO�O �O�O�O�O�O�O	__ -_?_Q_c_u_�_�_�_ �_�_�_�_oo)o;o Mo_oqo�o�o�o�o�o �o�o%7I[ m������ ��!�3�E�W�i�{� ������ÏՏ���� �/�A�S�e�w����� ����џ�����+� =�O�a�s��������� ͯ߯���'�9�K� ]�o���������ɿۿ ����#�5�G�Y�k� }Ϗϡϳ��������� ��1�C�U�g�yߋ� �߯���������	�� -�?�Q�c�u���� ����������)�;� M�_�q����������� ����%7I[ m������ �!3EWi{ �������/ ///A/S/e/w/�/�/ �/�/�/�/�/??+? =?O?a?s?�?�?�?�? �?�?�?OO'O9OKO ]OoO�O�O�O�O�O�O �O�O_#_5_G_Y_k_ }_�_�_�_�_�_�_�_ oo1oCoUogoyo�o �o�o�o�o�o�o	 -?Qcu��� ������)�;� M�_�q���������ˏ ݏ���%�7�I�[� m��������ǟٟ� ���!�3�E�W�i�{� ������ïկ���� �/�A�S�e�w����������ѹ�$FEA�T_DEMOIN�  ִ����ΰ�INDEX������ILE�COMP _w���7����-�SETUP2� `7�A���  N l�*�_�AP2BCK 1�a7�  �)�Ҹ�ϯ�%����ΰ :�����Ե��*߹�N� ��[߄�ߨ�7����� m���&�8���\��� ���!��E���i��� ���4���X�j���� �����S���w� ��B��f��s�+ �O����> P�t��9� ]���(/�L/� p/�//�/5/�/�/k/  ?�/$?6?�/Z?�/~? ?�?�?C?�?g?�?O �?2O�?VOhO�?�OO �O�OQO�OuO
_�O_ @_�Od_�O�_�_)_�_ M_�_�_�_o�_<oNo �_roo�o%o�o�oFɺz�P~� 2���*.VR�o�`* F�cLpZep�PCx��`FR6:��~\��{T��'��u�Q���x�w�Yf*.F
D���a	�s��Ռd�<����STM �"��-��p�Y��`i�Pendant �PanelY���H O���?���[�����GIF�6�A�"�ߟ8񟆯��JPG�����A���c�u�
��zJS��=��`У+��%�
JavaScrgipti���CSZ����@���k� %C�ascading� Style S�heets�_`
�ARGNAME.SDT�lD�\0Ϡ�P�`�q��`�DISP*g�J�D�����σ����ϡ�	PA�NEL1��O�%@D�8�x�k�}�+�2m߀��b���~ߐ�%�0�3 ��W�b�E����0�4u���b�����-��(�TPEINS.gXML4���:\H����Custom� Toolbar�����PASSWO�RD��}nFRS�:\���� %P�assword ?ConfigXo V��O��o�?� �u
�.@�d ��)�M�q �/�</�`/r// �/%/�/�/[/�//? �/�/J?�/n?�/g?�? 3?�?W?�?�?�?"O�? FOXO�?|OO�O/OAO �OeO�O�O�O0_�OT_ �Ox_�__�_=_�_�_ s_o�_,o�_�_bo�_ �ooo�oKo�ooo �o:�o^p�o� #�GY�}�� �H��l������1� ƏU������ ���D� ӏ�z�	���-���ԟ c������.���R�� v������;�Я_�q� ���*���#�`�﯄� �����I�޿m��� ��8�ǿ\������!� ��Eϯ���{�ߟ�4� F���j��ώߠ�/��� S���w߉���B��� ;�x���+�����a� ����,���P���t� ����9���]��� ��(��L^������� �$FIL�E_DGBCK �1a��� ��� ( ��)
SUMMA�RY.DG�h�MD:�0t �Diag Sum�mary1>

C?ONSLOG&	�t�CCon�sole log��=	TPACC�N�/%�4/?�TP Accou�ntin�>
F�R6:IPKDM�P.ZIPh/l
��/�/@P Exception�/n+�MEMCHECK�*/�@?�Me�mory Dat�aA?�LN�)	FTP��?'?�?�K7�mment� TBD�?u7 >�)ETHERNET�?f�!OHO�CEthern�et �figu�ra�/D�1DCSVRF�?�?�?�OQ1�%�@ verify all�OޗM,��EDI�FF�O�O�OO_R0{%�HdiffQ_�W�!�@CHGD1pF_-_?_�_ f_,�_S+P�Y2�_�_�_Xo �_oo�GD3No5oGo�o� no�fUP?DATES."p~iFRS:\ �a}DUpdates Lista�fPSRBWLD'.CM�hLr��c�PS_ROBOOWEL�?<�aHADOW�o�o�o�f�Q3Shado�w Changeysi��=�&�NOTI�OA�S���O5Notifi�cqB���O�A J?�nc��p���D ��L��󟂟���;� M�ܟq� �����6�˯ Z��~���%���I�د m�����2�ǿٿh� ����!�3�¿W��{� 
ψϱ�@���d���� ��/߾�S�e��ω�� �߿�N���r���� =���a��߅��&�� J���������9�K� ��o����"�����X� ��|�#��G��k }�0��f� ��,U�y ��>�b�	/� -/�Q/c/��//�/ :/�/�/p/?�/)?;? �/_?�/�?�?$?�?H? �?�?~?O�?7O�?DO mO�?�O O�O�OVO�O zO_!_�OE_�Oi_{_�$FILE_Lp{PR[p��_P����X�MDONLY 1�a�UZP 
 �
_�_._oR_o;o __o�_�o�o$o�oHo �o�o~o�o7I�o m�o� ��V� z�!��E��i�{� 
���.�ÏՏd����� ���*�S��w���� ��<�џ`������+� ��O�a�🅯���8����߯�ZVISBC�K�X�Q�S*.V�D�0���FR:�\��ION\DA�TA\�â���Vision V?D file\�j� ����̯ڿį����� 4�ÿX��|ώ�ϲ� A���e�w�ߛ�0�B� ��f��ϊ�ߛ���O� ��s����>���b� ����'������� �����'�L���p��� ����5���Y���}����$�ZMR2_GR�P 1b�[��C4  B� 	� �Qk}h E��� E�  F?@ F�5U�/
�h L���M���Jk�K�v��H�,�Hk�=�?�  �/�h 9tQv8�?��6h�%��A�  3EBH�eB�a `�E@�i/g��h @�UUU�U��>�]�>П��;r8	==�=E��<D�>�<�ɳ<�Ε��:�b�:/'�79�W�9
@��8�8�9���T/�Q/�/eE�7� E?p D�D�/�D�  ?D�  Cζ/9
_CFG c�[T �/?0?B?��NO �Z�
F0x1 }0�R�M_CHKTYP  �P� �P�PڟP��1OM�0_MsIN�0
���0v�PX�PSSB�#]d�U�Pi��?	�3O$O�UTP_DEF_OW�P�
�Y?AIRCO�M�0JO�$GENOVRD_DO�6��RxLTHR�6 �d�Ed}D_ENB�iO }@RAVCrGe�7� ���FnH E�� �Ga H�� �H�@Jh`�/O?_�G_X_{� ��AOU�@kN {NB{8���_y_�_��_�_  C�� 	�$o�XYoilCOmB���AVb~	�Y+O�@SM�T�Cl�IZ �04d��$HOSTC�"1�m�� 5	
x
{
:byeV�� ���zu� ��$��GH��p	anonymousK�y��� ������	-� A�c�V�h�z���� ��ԟ����M�_� @�R�d�v���ˏݏ� ���7��*�<�N� `�����������̿� !�3��&�8�J�\ϟ� ��ïկ׿������� �"�4�w�X�j�|ߎ� ������������� 0�sυϗϩϫߜ��� ���������K�,�>� P�b���s��ߪ����� ����G�Y�k�L� p�������  $6YZ��~ ����	�-?  /SuB/h/z/�/�/ ��/�/�/�/
?-/_ qR?d?v?�?�?�� //?�?I/*O<ONO `OrO�/�O�O�O�O�O O3?E?&_8_J_\_n_��g�aENT 1n~�i�  P!�O.�_  �@�_�_ �_o�_+o�_Ooo[o 6o�o�olo�o�o�o�o �o9�oo2� V�z����� 5��Y��}�@�v��� ��׏��������+� �T�y�<���`����� 埨�	�̟ޟ?��c��&���J�QUIC�C0��p�!17�2.8.9.22	5����1�����3�¦�24��"���!?ROUTER��`��r�ӿ!PCJO�GԿ��!19�2.168.0.�10����CAMP�RT$� �!�1�K�2�RT��O�a���ψTNAME �!�Z!ROBO�=���S_CFG �1m�Y ��Auto-s�tarted�4FTP�?[��?�O ��O�߼������ߋO �(�:�L�o�]��� ���������04�F� X�9�l��P������� ��z�������#F� ��Yk}����?�=SM�65233)�
=_�,R dv�K���� �ӯ�3/E/W/i/{/ $q��?�?�? �/3?&?8?J?\? /�?�?�?�?�?�/m? �?O"O4OFOXO�/�/ �/�/�?�O?�O�O_ _0_�?T_f_x_�_�_ �OA_�_�_�_oo,o oO�O�OEo�_�o�O�o �o�o�o�o(:L ^�o����� � �CoUogoH�{�o �������Ə���� � �2�U�׏U�z��� ������)�;�� O�q�R�d�v�����]� ��Я����)���<��N�`�r�������_ERR o�ʡ����PDUSIZ  �3�^L��ȴ>~�WRD ?"����  guest-�!�3��E�W�i�{���SCD�MNGRP 2p�"�˰���3��-�K�� 	�P01.05 �8�� �����>� j  2�1��� � ����T��������������$Ё��ϿQ�<�u�`�������  ��  
���N(�P,�(�����Q����������l�� 8�#{�d�����"ߙ�__GROU��q�������	����4�S�QUPD  d�ȵX��TY������TTP_AUTH 1r��� <!iPeOndan����8��g�!KARE�L:*����K�C-�=�O�%�VI�SION SETb�����!������ "� ��_6H�l~��CTRL s�����3����FFF9E3���FRS:D�EFAULT�FANUC W�eb Server����	�Ĵ}��������WR�_CONFIG ;t�� ���IDL_CPU_kPC*3�B���I  BH/%MIN�:,��M%GNR_I�O�����Ƿ1 NP�T_SIM_DO�&�+STAL_oSCRN& ��*�TPMODNTOqL�'�+bRTY�(pI!�&����ENB�'���-$OLNK 1u���Q?c?u?��?�?�?�?52MAS�TE~ ��52SLAVE v��34��O_CFG�?IU�O��OBCYCL�E>OD$_ASG� 1w����
  �?�O�O�O�O�O�O_ _1_C_U_g_y_�_�;�tBNUM�Ĺ
BIPCH[O��@RTRY_CN*��"ĺB�!���P1�bȵ B;@Bx�>��Jo�1 SDT_ISOLC  ���f��$J23_�DS4�:��`O�BPROC?�%J�OG^�1y�;���d8�?���[�o�_?؟֟O|Q Ns��V����-�~o�h�`Y A|�_�bPOSRE�o~�&KANJI_�0����/k�+�MON #zg��2�y�Ϗ�����Ҿ)�0c{�,�9�T���e�_�LY �R�_k�EYL_OGGIN@�����ȵ�$LA�NGUAGE ,k2$ 㑱��LG1b|�2���R3�x������O �� '0,�� կ
q�3�M�C:\RSCH\�00\��LN_DISP }�?bf�MKm�OC�"�@"Dzh#�A�O�GBOOK ~�K��w���w�w���X���-�?�Q�c�u�`��11����	� ��h�޿����ॐ�_BUFF 1@=���)��� ��E�a�sϠϗϩ� ���������B�9� K�]�oߜߓߥ��ߜ�~�DCS �� =��͗�ֿM��l:�L�^�p���IOw 1�K No������������� ��%�9�I�[�m��� ���������������!3EY��Ex TMlnd����� �0BTfx �������/8/���SEV`}�]�TYPln�`�/�/�/)-P�RS�P����bFL 1���`��?,?>?`P?b?t?�?�/TP���loq"��NGNA�M�d��Ւ��UPSFu�GI�U\�e�1�_LOAD�`G {%}�%DF@�GI6�?�[MAXUALRM�Wk�X�\@�1_PR�T`hԣ��Z@Cx�������OV�9ŜC�`P �2��K �9�	�q!P]  ��OQ�R9_$_6_o_ �]_�_�_�_�_�_�_ �_oo@oRo5ovoao �o}o�o�o�o�o�o *N9rUg� ������&�� J�-�?���k�����ȏ ڏ�����"���X� C�|�g�������֟�� ��ݟ�0��T�?�x� ��m�����ү��ǯ� �,��P�b�E���q����SGD_LDXD�ISA�0�;��ME�MO_AP�0E {?�;
 j  ����*�<�N�`�r����Z@ISC 1��; �����T�A����ϛ�$��Hߙ�C�_MSTR ��B-g�SCD 1����<߶�8������� ��"���X�C�|�g� ������������� 	�B�-�f�Q���u��� ����������, <bM�q��� ����(L7 p[����� �/�6/!/Z/E/W/ �/{/�/�/�/�/�/�/ ?2??V?A?z?e?�?��?�?X�MKCFG� �vݽO�CLT�ARM_�2��G�B P�2�@>OFD{@�METPU�C�@��~�ND�@ADC�OL`E�@kNCMN�T�O tEo� �v��N5C.A�O�DtE_POSCF�G�N�PRPM�OYST�@1��� 4@��<#�
oQ�1oU _�Wk_�_�_�_�_�_ �_o�_oOo1oCo�o goyo�o�o�o�o�atA�SING_CHK�  �O$MODAQC��?���>+u�DEV 	��	�MC:_|HSI�ZEѽ���+uTA�SK %��%$�12345678�9 ��u)wTRI�G 1���l#E% ��)����S�6�%C�v�YP�q>�At*sE�M_INF 1��#G `�)AT&FV0�E0`�׍)��E�0V1&A3&B�1&D2&S0&�C1S0=ƍ)GATZ׏+��H/� W��K���A���� j�ӟ����	� ��.� ������;���� Я⯕����*�<�#� `��%���I�[�m�޿ 鯣��K�8����n� )ϒ�y϶���{��ϟ� ��ÿտF���jߡ�{� ��S����������� ����T���+ߜ�� a���	�����,��� P�7�t���9��]�o� �����(:q�^ ��=����X�NITOR�@G �?s{   	�EXEC1�32*%3%4%5%�p�'7%8%9�3  ��$�0�< �H�T�`�l��x���2�2��2�2�2�2��2�2�2�2*�3�3�30+q�R_GRP_SVw 1��� (�a���:��hK�=�&7��);��=>�T�E�av�q_D{�~�1P�L_NAME �!#E0�!D�efault P�ersonali�ty (from� FD) �4RR�2�! 1�L6�8L@�1P
d d�?v?�?�?�? �?�?�?�?OO*O<O NO`OrO�O�O�O�O�O�OJx2e?_ _2_D_�V_h_z_�_�_�_r< �O�_�_�_o"o4oFo�Xojo|o�o�o�i�VD�_�n
�o�oNtP�o *<N`r��� ������&�8� n���������ȏ ڏ����"�4�F�X� j�|�K�]���ğ֟� ����0�B�T�f�x����������Ү �FnH F�� �G=��'�   �����"d���0� B�&�d�r��׭Ҫ\�੿����ݿ�  ͸��� ��0�6�T��vϿ �ϩ�ͰA�  ��˿��Ǹ]0 ���ƿ3�¿W�B�{� ��x߱�B5K3�9^0�`�!0 �� �0�� @D7�  ��?�����?� ��!A������$��(;�	l��	 ��p�V� ]0M�� � � � ��l�r� K(���K(�K ���J�n�J�^/J&Ǔ�2�������� @Y�,@�Cz@I�@��������N�ߠ��f���_��I���S�z��Ä��  <���% �3�������!?s8y�
��/�!�x����T� ܌���������}��  _  �����o�  ����������	'� �� 0I� ��  �����:��ÈTÈ=�c��l��	�(|@�����Ѧ�������N@0�  '�� ���@2�@���@!�����@)��C@0C�W�\CI�CM�CQ��� ��ģ��%%���/� ��B���@0��l@� ��!Dz���V�//+/�Q/���� �aH@q)q�%  �S�+��� p�!?�ff���/�/V/C ���/;��8�  !?/:��D4�� \6�Pf8�)c�\�\��?�Lv �$��;�Cd�;�pf<߈�<��.<p��G<�?L:��ݧA����d����?f7ff?�?&@���@�� B�N�@T�,E�	��	A ���dO�O�7H� �/�O�O�O�O _�O$_�_H_Z_E_~_�MEF�m_�_i_�_UO�_�yI�_2o�XC��E���"Gd G; ML!o�omo�o�o�o�o �o�o�o$H��i ww9��_�o�U ��*�<�ڪ����/ �6������ď���
��A�A������C؏=�ԏ��X���񨑟,�����  ģP��"@�<��E� C���s��x��؄�(�����/�B��/B"�}A���#A��9@��dZ?vȴ,���~��<)�+� =�G���j���q���
�AC
=C������년� ���p�Cc�����B=���ff�{,��I���HD-��H�d@I�^�?F8$ D;ޓܪ��̠Jj��I��G�F�P<���QpJn�PH�?�I��q�F.� D� �Ɵg�R���v����� ���п	���-��Q� <�Nχ�rϫϖ��Ϻ� �����)��M�8�q� \ߕ߀߹ߤ߶����� ���7�"�[�F�k�� |�����������!� ��W�B�{�f����� ����������A ,eP�t��� ���+;a�L�p�����(�����3:��1�y�%�3�V��/"�(/:/�!�4M��T/f/F1��=Ӏ/�/4Ue'��T9�-�)�/@�/?�/4?"<]�P�2	Pf>�q��?��?��?�?�?�9���( �?�?/OO?OeOPO�QB�hOzO�O�O�O�O��O�?t.__R_@[/X_b_�_�_�_�_�_�Q{f�_�_o
o@o�.odorj  2 wFnH"�F��"��G=��B# ��C9)��@|�@��o ��q�o{E�� F}��`�H C������oA`��kE�0wGa�O����{Q?ސ�q �\d � zq `�
 �!�3�E�W�i� {�������ÏՏ��������q ��P+��~Y��$MSK�CFMAP  ��%� �^f�q�qp�D�ONR�EL  X5�[��0D�EXCFE�NB��
Y����F�NC����JOGO/VLIM��d����]dD�KEY����=�_PAN���\�D�RUN����>�SFSPDTY�w0������SIGN|����T1MOT����D�_CE_G�RP 1��%[�\�O��O�&��d �Q��u�,�j���b� Ͽ��Ŀϼ�)�;�� _�σϕ�LϹ�pϲ� �Ϧ��%��I� �m���fߣ�OvD�QZ_�EDIT��U��T�COM_CFG 1�Q�����"�}
��_ARC_���X5ؙT_MN_oMODE��縙UAP_CPLF����NOCHECK� ?Q�  W5�H���������� '�9�K�]�o������������v�NO_WA�IT_L���׾�NMT���Q��{o_ERRȡ2�Q��1� ��t����H*�����`�O�I�Px b<���!8�?�0|4�pBPA�RAMJ�Q����	��7so� �=�`345678901�/ *�?/ Q/-/]/�/�/u/�/�/�+�7�?<�7?���UM_RSPA�CEN�'2$�p?z4�$ODRDSPE������OFFSET�_CAR�Ќ�6D�IS�?�2PEN_FILE�0�$�����1PTION_I�O
�=�@M_PR�G %\:%$*�IO[N�3WORK ��Χ�� ����F7��Bh�� ɢ�d�@(7�A	 a��x�A5��c��0�RG_DSBL  \5���|_�1RIENTTO��9�C��pZ��a�0�UT_SIM_D�GX�+��0V�0LCT �%�ҟD<x=gT_PEXh��?n�TRATh� d����T�0UP �u^�Ӡ�oo�_�:oHi�$�2ǣ��L68L@�>_S
d d'?�o �o�o�o�o�o�o 1CUgy��� ����I2~o'� 9�K�]�o���������ɏ9�<����)� ;�M�_�q��������� H�j3�H1`��XRP�C�U�g�y��� ������ӯ���	�� -�?�Q� �2������� ��Ͽ����)�;� M�_�qσϕ�d�v��� ������%�7�I�[� m�ߑߣߵ�����X�ϡ��*��S�H�Z�?�}������ &?��������� ���+�I�O�m�����?@����� A�  �������� ��M8q\�����z�d`O�P1��k����sd`�R0 ���D$@ @D� � DD?QD�	��U�  �;�	l1	 ���p��s& ' j � �/ � ʉ�� �H<zH<W��H3k7G�CG���G9|+c�	�H
��� CC
9P/9P49S;Q9/���9  �� � 1!�H7 3�����/1/C/�BY�����XQ��^�H�<Pq/ ܀�/�"2�#�3�.��    ��0�� �  �0�6�/?�	�'� � M2�I� �  y���
=���q?�;�#&�(�3�/��A�?4;�B�?�9NEPO  'VP3D��b CEPC��\Cf Cj Cn/@ORO>ߑ  ����D�%%�_�� �B��0�FEP�E˜@XP�E5z�_s/8_#_H_�n_�"�� �aH]2�Y�A�U  �CS�H�A�0p�Q?�ff���_�_s_C ��o(k�18�0 >oLj-�!adTW�0yf�P�h�Y�yy�3?�L�0�T�!;�Cd�;�pf<߈�<��.<p��G<�?ij��WA�E�ل1d�31��?f7ff?�@?&+pVT�@��=r�N�@T�IuՉ��&q -�0!��we  o������A� ,�e�w�b�������я ����l���O���CE���2Gd G;�|>����� ß���ҟ����A� ,�e�����V���� د6���r�#�5�G�Y��Z� �_�f��������̿��A @A�@%���5�C��Z��<�/i�?�؈Ϗ�8�ϳ�U�P��2]!zYNE� CU�%�̣�Ŀ����E�@�I�!t�B�/�B"�}A��#�A��9@�dZ�?vȖ+~��~�����<)�+�� =�G�(߇Ԁ��q���
AC�
=C������녡� ��p��Cc�¥��B=���f�f�{��I����HD-�H��d@I�^�F8�$ D;���ڭ���Jj��I���G�FP<���QpJnP�H�?�I�q�?F.� D��E�� ��o��������� ��&��J�5�n�Y�k� ��������������  F1jU�y� �����0 T?xc���� ���//>/)/;/ t/_/�/�/�/�/�/�/ �/??:?%?^?I?�? m?�?�?�?�?�? O�? $OOHO3OXO~OiO�O��O�O�O�O��(}��g�3:�O�a��)U�E3�V�_+_9R��E_W_t�4M㇬q_�_t��=�ӝ_�_4Ue'��T9�]�Y	o�_-oPoQo?lz�P�bP�n�����o�O�o�o�o<�i���(�L7\�mt�B� ��������o`��K�9�o�]�/u�������ŏ�ُ�{f��9�'�]�K������  2 Fn�H��F�Щ�G=b��B@P!�.�C9F��p��@2���	��C��E�� F����H C���S�b����������¯ԯ���?����y�RC�C�|�C�}�
 ۯ>�P�b�t� ��������ο���p�(ϧ�� ��m[��~Y��$PA�RAM_MENU� ?�U��  DEFPULSE4��	WAITTM�OUT��RCV��� SHEL�L_WRK.$CUR_STYL��;��OPT��ϧPTB����C��R?_DECSN��te G�A�S�eߎ߉ߛ߭� ����������+�=��f�a�SSREL_�ID  �U�a��u�USE_PRO/G %p�%b���v�CCR����ax����_HOST �!p�!�����T �`��8����:�t�>��_TIME�����a�GDEBU�G��p�v�GINP?_FLMSK����sTR����PGA��e ��{�CH��^��TYPEm�y�a�[����� �!JEWi �������� "////A/j/e/w/�/ �/�/�/�/�/�/??�B?��WORD ?�	p�
 	RyS��	�PNSu���~2JO�
��TE[��?COL�u>8�?>L�� ��P��p���TRA�CECTL 1�v�Uz� �`L ������1L�FDT Q��U�^@#@D � nsc/3BkO}I{O�O�D��O �O�O�O�O_%___ []�Oe_�_9_�_�_�_ �_{_�^o�_�_Tofo xo*o<o�j�o�o�o�o /ASew� �������� +�=�O�a�s������� ��͏ߏ���'�9� K�]�o���������ɟ ۟����#�5�G�Y�k�}���gI���� ӯ���	��-�?�Q� c�u���������Ͽ� ���)�;�M�_�q� �ϕϧϹ�������� �%�7�I�[�m�ߑ� �ߵ����������!� 3�E�W�i�{���� ����������/�A� S�e�w����������� ����+=Oa s�������� '9K]o� �������/ #/5/G/Y/k/}/�/�/ �/�/�/�/�/??1? C?U?g?y?�?�?�?�? �?�?�?	OO-O?OQO cOuO�O�O�O�O�O�O �O__)_;_M___q_ �_�_�_�_�_�_�_o o%o7oIo[omoo�o �o�o�o�o�o�o� EWi{��� ������/�A� S�e�w���������я �����+�=�O�a� s���������͟ߟ� ��'�9�K�]�o��� ������ɯۯ���� #�5�G�Y�k�}����� ��ſ׿�����1� C�U�g�yϋϝϯ��� ������	��-�?�Q��c��$PGTRA�CELEN  �b�  ���a��w�_UP �����љ�В���w�_�CFG ������a���������������aл�DEFSPD ����`щ��w�IN~��TRL ������8�F�PE_C�ONFI�Ш��O������WLID�ө��	��LLB 1���� t�?B�  B4��� ��� ����� 88�?�0�K�0�G�i�k�}� ������������5Ak��� ��2��	�?~��GRP 1����lb�A�  ��333a�A���D�@ D�� �D@ A@�Ta�d+������� 	='����#´#��B 9!�///O/9/s/
?��?����/�/��.�/ =o=	7L�/?�/?P? ;?t?_?�/�?�??�?<�?�?  DzC Oa�
OHO�?XO~OiO �O�O�O�O�O�O_�O�_D_/_h_S_�_�Z!�a�
V7.10�beta1�� �Ax���R�y�y�Q?���Qo>�\)�QB0����PA��SBp���QA�9Sy�b
a�S �_2oDoVoho��Ap���"���o��o�o�o�Ҹө�KNOW_M  �|�֦�SV ���/���5O8 J\u_�k}��Ҕ���M]�z�Д��R	��a�%%��"��|���� ��u��P@ �a�]�a�q�m��`��MR]��}��&%O`�P�$ӏ�KST]�1 1���
 4��vi�Q:��"�4� F�w�j�|�������ğ 	����?��0�u�T� f����������ү���2� �a��<K��^35�G�Y�k��4���������A5ۿ�����6.�@�R�d��7�ϓϥ����8������
���MAD  �����OVLD  ���G�PARNUM  ��|����T_SCHy� ��
�����0�UPD��������_CMP_�p|�p�p'�e��ER_wCHK�����j����RS��oWG_MO{���_��~��_RES_G��� o��������� ������2%V�Izm`�R�4�\� l��Q������S� ڰ�S�-�9X ]S��x��S��� ���S�&��//S�V 1���a�q�@c?\�THR_INR��~��rz�ed�&MASS�/� Z�'MN�/�#M�ON_QUEUE� ���f"��a*��N��U��N�&��0END1;�79EcXEF?75\�BEE0|'?3OPTIO$7�D�0PROGRAoM %�*%0�T/��2TASK_�I{ԍ>OCFG ���/���?"@DAkTA�s�+K��"�2��O�O�O�O�O �O�O_!_3_E_�Oi_�{_�_�_ROINFO
�s�oM�
4[_�_
o o.o@oRodovo�o�o �o�o�o�o�o*�<N`�W�T�oL ��	!A�K_%Aq�+I�^�vENB|�H�})��v2��xG%A�2��{ P(qO�4�F� C��e��z_EDIT ��+O����DWE�RFLg8|# �RG�ADJ ��:A	����?"���!߆�1�q�]�g�?���A<@��v%<�l�ӈ���q�2�)��R	H0l�e�{"6�?
���AF$�t$ܖ�*�/� **: ��"�����d�1�f�Ցd�[�_"U�#��� 3�E�s�i�{������� ߯կ�a���K�A� S�Ϳw���������9� ���#��+ϥ�O�a� �υϗ�߻������� �}�'�9�g�]�o��� �ߥ�������U���� ?�5�G���k�}��� ��-���������� C�U���y������� ������q-[Q c������I �3);�_q���t&	>O@/Հ ./g/R$ݙ�/ߓU/�/�Q/�/�/�PREF� �)�ՀՀ
~߅IORITY�7�2F��MPDSP�1яG7UTFǓކ�ODUCT
A��:�/��OG��_�TG΀B���2TO�ENT 1�� (!AF_I�NEq0OG!�tcpO6M!�ud%O^N!iccmMOu��2XY"��Í��X1)� 0��O�OX0��O�O �E�O)__M_4_F_�_ j_�_�_�_�_�_o�_$%o7o*�3"��=Y�xyo�o��>��J���/�io�o���􂘅�AK�,  �0�q'9K]�X5�7�pHANCE� �)��rrn{d �o��uyw	3�?"3�ق�PORT_N�UMr3X0����_CARTRE�PR0����SKST�Aq7 C�LGS6 @ȍ��K�X0�Unothing�����̏܌������#��?k�TEMPG ɕ94�����_a_seiban�/���/��͟��� ܟ� �9�$�]�H�Z� ��~�����ۯƯ��� �5� �Y�D�}�h��� ��ſ��¿����
� C�.�g�R�wϝψ��� ������	���-��*� c�N߇�r߫ߖ��ߺ� �����)��M�8�q��\��6�k�VERS�IP0�7�� disable�r�<�SAVE ���:	2600H�844����,�!`�.�@�_Od� 	��H{2 /����X�e�� ��	-;
��c��n ��L��_�0 +1˧K�� "�����0URG�E�pB�0T6>5�W�F� DOr6�r�6W��0�"�WRUP�_DELAY ��;�R_HOT %%&~1��+�R_NORMAL�y�2���SEM�I��"/�!QSKKIP���w�x�� g/��/�/�/r-�5�/ �'�/??(?�/L?:? \?�?�?�?l?�?�?�?  OO�?"OHO6OlO~O �OVO�O�O�O�O�O_ �O2_ _V_h_z_@_�_��_�_�_�_�_���$�RBTIF?�R�CVTMOUT�vB��`DCR�}�E) �~!�7���C����C���A7�f��/|#�lD��i���$�a9r/��o�o ;�Cd�;�pf<߈�<��.>�]�>П��o��o'8} 8^p� ������ ���$�1%RDIO_T?YPE  ��.�EFPOS1 �1���  x �����Ώ���{� ���:�Տ7�p���� /���S�ܟ���՟ 6�!�Z���~����=� ��دs����� ���D� V���=�����¿]� 濁�
ϥ��@�ۿd� ����#ϬϾ�Y�kϥ� ���*���N���r�� oߨ�C���g��ߋ�� &������n�Y��-� ��Q���u������4� ��X���|���)�;�u� ����������B�� ?x�7�[� ����>)b� �!�E��{/ �(/�L/^/�/E/ �/�/�/e/�/�/?�/ ?H?�/l??�?+?�? �?a?s?�?O�?2O�? VO�?zOOwO�OKO�O oO�O�O_._�O�O_ v_a_�_5_�_Y_�_}_ �_o�_<o�_`o�_�o<�o|�2 1ш�2o Do~o�o�o &oD�o he�9�]� �
�����d�O� ��#���G�Џk�͏� ��*�ŏN��r��� 1�k�̟��🋟��� 8�ӟ5�n�	���-��� Q�گu�����ӯ4�� X��|����;���ֿ q�����Ϲ�B�ݿ� �;Ϝχ���[���� ߣ��>���b��φ� !ߪ�E�W�iߣ���� (���L���p��m�� A���e�������� ���l�W���+���O� ��s�����2��V ��z'9s�� ���@�=v �5�Y�}� ��</'/`/��// �/C/�/�/y/?�/&? �/J?�/�/	?C?�?�? �?c?�?�?O�?OFO �?jOO�O)O�O�o�d3 1ҵo_OqO�O )__M_SOq__�_0_ �_�_f_�_�_o�_7o �_�_�_0o�o|o�oPo �oto�o�o�o3�oW �o{�:L^� ����A��e� � b���6���Z��~�� ����Ə �a�L��� � ��D�͟h�ʟ���'� K��o�
��.�h� ɯ�������5�Я 2�k����*���N�׿ r�����п1��U�� y�ϝ�8Ϛ���n��� ��߶�?�������8� �߄߽�X���|��� �;���_��߃��� B�T�f�����%��� I���m��j���>��� b����������� iT�(�L�p ��/�S�w $6p���� /�=/�:/s//�/�2/�/V/�/�O�D4 1��O�/�/�/V?A? z?�/�?9?�?]?�?�? �?O�?@O�?dO�?O #O]O�O�O�O}O_�O *_�O'_`_�O�__�_ C_�_g_y_�_�_&oo Jo�_no	o�o-o�o�o co�o�o�o4�o�o �o-�y�M�q ���0��T��x� ���7�I�[������ ���>�ُb���_��� 3���W���{������ ß��^�I������A� ʯe�ǯ ���$���H� �l���+�e�ƿ�� 꿅�ϩ�2�Ϳ/�h� ό�'ϰ�K���oρ� ����.��R���v�� ��5ߗ���k��ߏ�� ��<�������5��� ��U���y������8� ��\�������?�Q� c�������"��F�� jg�;�_����/45 1� ?���n�� �f���%/�I/ �m//�/,/>/P/�/ �/�/?�/3?�/W?�/ T?�?(?�?L?�?p?�? �?�?�?�?SO>OwOO �O6O�OZO�O�O�O_ �O=_�Oa_�O_ _Z_ �_�_�_z_o�_'o�_ $o]o�_�oo�o@o�o dovo�o�o#G�o k�*��`� ���1����*� ��v���J�ӏn����� �-�ȏQ��u���� 4�F�X����ޟ��� ;�֟_���\���0��� T�ݯx���������� [�F�����>�ǿb� Ŀ����!ϼ�E��i� ��(�b��Ϯ��ς� ߦ�/���,�e� ߉� $߭�H���l�~ߐ��� +��O���s���2� ����h�������9�<16 1�<�� ��2������������� ��R��v� 5�Yk}� <�`���� U�y/�&/�� �/�/k/�/?/�/c/ �/�/�/"?�/F?�/j? ?�?)?;?M?�?�?�? O�?0O�?TO�?QO�O %O�OIO�OmO�O�O�O �O�OP_;_t__�_3_ �_W_�_�_�_o�_:o �_^o�_ooWo�o�o �owo �o$�o!Z �o~�=�as �� ��D��h�� ��'���]�揁�
� ��.�ɏۏ�'���s� ��G�Пk������*� şN��r����1�C� U����ۯ���8�ӯ \���Y���-���Q�ڿ u�����������X�C� |�Ϡ�;���_����� ��߹�B���f�L�^�7 1�i��%�_� ������%���I��� F����>���b��� ������E�0�i�� ��(���L������� ��/��S�� L ���l��� O�s�2� Vhz�/ /9/� ]/��//~/�/R/�/ v/�/�/#?�/�/�/? }?h?�?<?�?`?�?�? �?O�?CO�?gOO�O &O8OJO�O�O�O	_�O -_�OQ_�ON_�_"_�_ F_�_j_�_�_�_�_�_ Mo8oqoo�o0o�oTo �o�o�o�o7�o[ �oT���t ��!���W��{� ���:�Ï^�p����� ��A�܏e� ���$� ����Z��~����+� Ɵ؟�$���p���D� ͯh�񯌯�'�¯K���o�
���yߋ�8 1ז�@�R���
��� .�4�R��v��sϬ� G���k��Ϗ�߳��� ���r�]ߖ�1ߺ�U� ��y�����8���\� �߀��-�?�y����� ���"���F���C�|� ���;���_������� ����B-f�% �I���, �P��I�� �i��/�/L/ �p//�///�/S/e/ w/�/?�/6?�/Z?�/ ~??{?�?O?�?s?�? �? O�?�?�?OzOeO �O9O�O]O�O�O�O_ �O@_�Od_�O�_#_5_ G_�_�_�_o�_*o�_ No�_Ko�oo�oCo�o go�o�o�o�o�oJ5 n	�-�Q�� ���4��X��� �Q�����֏q����� ����T��x�����7�������MASKW 1�û������XNO  ����MOTE � 3����i�_CFOG �p�����PL_RANGl��g�t�POWER ��õݠ|�SM�_DRYPRG �%p�%m���T?ART �ծ#�UME_PRO������_EXEC_ENB  d�=x�GSPDX���v����TDB���ϺRM޿ϸI_A�IRPUR�� pp�B�<�ٛMT_��TРn��OBOT_ISOLC1���8�����9�z�N�AME p��n�ۙOB_ORD_NUM ?ը�5�H84�4 g��b�Ҙ ����/(/�^/�Ҧ/���PC�_TIMEOUT��� x�S232扢1�4�γ L�TEACH ?PENDANPЅ�,������l�j��Mainten�ance Con%sg��߾�"��f�No Use�� �߮���0�B�T�⒎h�NPO2�RҤ��z�e�CH_�L[��p���	����!UD1:����R�VAIL���R����x�e�PACE1 2�p�
 �濫��{鈋�������9˺�8�?�%���%� ��4IDu��� ����Y������ ):!4�8�Uu� �����/� ):/!/O/q��� U/���/ ?�/?6? ?K?m//�/�/�/c? �/�/�/�?O2O	OO i?{?�?�?�?_O�?�? �OGO_._@_'_eOwO �O�O�O[_�O�O�_o �_+_<o#oQos_�_�_ �_Wo�_�_�o�o 8Moo�o�o�o�o �o�o�D��4�� I�k}���a�� �돽��0�B��+�
X�2a�s������� W�͏�����4�U�<�j�o�3~������� Ɵt����<���Q�r�Y���o�4������ ѯ㯑��)�8�Y�� nϏ�vϤ�o�5��ʿ ܿ� Ϯ�$�F�U�v�@9ߋ߬ߓ���o�6�� ��������A�c�r�V�������o�7 ����(�:���^�� ����s���������o�8�!�3�E�W�{� ��������o�G �/� m�
u d  /���� ��/Nl -S-L/�/p�d� z� �/�/�/�/??&?/ ./@.1:n?�;�?�/�/ (?�?�?OO*O<O2? D?V?h?�?�O�O�?�? HO__&_8_J_\_RO�dOvO�O�O�_ ` @p��U]/o�O�IAakU�_Rodo j_DjEowo�o�o�o�o �o%�o�o= ASe���	�� �3�E���+�]����a�o\
#o�o�_M?ODE  /
�/S �/㏙_��Z�oH�����	���㟐�CWORK�_AD�
��@^��R  /< �1���_INTV�AL�a�%�R_�OPTIONR� �%���V_DA�TA_GRP 2Y�uX:D�@PП ��̟�˩͏���1� �U�C�y�g������� ӿ������	�?�-� O�u�cϙχϽϫ��� �������;�)�_�M� ��qߧߕ߷������ ��%��I�7�Y�[�m� ������������� �E�3�i�W���{��� ����������/ SAwe�����P�$SAF_D?O_PULS�Q�A��� CAN_GTIM��E}��R ���Ƙ_qsy�֡��Yo�K�C կ������ l//%/7/I/[/e�+�C�2�$K�)d�$�!ѢIf)�P5��/�/�/���)��/ ��4�_; �R  T0�!?�^?p?�?�9T D���?�?�?�?�? O O$O6OHOZOlO~O�O��O�O�O�OU�s��'��O$_6_�I � �T;�o���WQo�p�M
�t��Di��[=Z?0 � ��o� [Q[SC�_�_�_�_ o o2oDoVohozo�o �o�o�o�o�o�o
 .@Rdv��� ������*�<�@N�`�r��������? ��я�����+�=� O���r%{�������ß ՟�����"�_���02�SwU�]n����� ����ȯگ����"� 4�F�X�j�|������� Ŀֿ�����0�B� T�f�xϊϜϮ����� ������,�>ߩ�b� t߆ߘߪ߼������� �o�(�:�L�^�p�� ����#�Q�[���� 
��.�@�R�d�v��� ������������ '9K]o��� �����#5 GYk}�������O�3�// 1/C/U/g/y/�/�/�/ �/�/�/�/	??-?;:��D?q?{6���d�j?@]	12�345678�R�h!B!��*��B��V��? �?OO)O;OMO_OqO wA��O�O�O�O�O�O __*_<_N_`_r_�_ �_�_�_�]�O�_ oo $o6oHoZolo~o�o�o �o�o�o�o�o�_�_ DVhz���� ���
��.�@�R� d�#��������Џ� ���*�<�N�`�r� ��������y�ޟ�� �&�8�J�\�n����� ����ȯگ����ϟ 4�F�X�j�|������� Ŀֿ�����0�B� T�f�%��ϜϮ����� ������,�>�P�b� t߆ߘߪ߼�{����� ��(�:�L�^�p�� ���������� ����0.�@�%���l��~����Cz  �B\�   ���2d4� ���d1
���  	�d22,�%7,IXp���Z������� %7I[m� �������!/ 3/E/W/i/{/�/�/�/ �/�/�/�/??/?A? S?e?w?�?�:Z������<�4��`�$S�CR_GRP 1��� ��� �� ���� ��	 /�1��2
B D[����� I�7GDO82OkO�����hBDE� DP�w�C�GhK�AR�C Mate 1�20iC 678�90��M-�@A� 8��M2IA��A��
1234�5�D;F�2  ����>U�1{F�1HC�1�AhAJ<ANY	?R�_�_�_�_�_�\?��H��0�T�7�2 o/O0oVoho7F/��Co�o?o�o`���l0Q�o:DBǲ�!�r2tAA��A�  @��YuA@��Wpj ?�wrH��DzAF@ F�`�r��o�� ���B�-�f�Q��� }Yq�r������ďքB��y�*��N�9� r�]�o�����̟��� ۟�&���CTOF�k�����h�����qYqO6���7G@Yp4ݯ����W\HC+�3���AnpC�V�$�o~ec��W���A y���������ո���¿ P�(��%�7�I�v�b�SS���0EL_DEFA�ULT  m�����u�HOTSTR�͐����MIPOWERFOL  ������oWFDO�� ��� u�RVENT �1���`��� L!DUM_�EIPL�(��j!AF_INE��<Fߺ�!FT�u��<ߙ�!o�� ������!RPC�_MAIN���غ8��1���VIS���y� �}�!TPp��PUt�/�dl���!�
PMON_PR'OXY��2�e���Ȑ���+�f�a�!RDM_SRVb�r/�gP���!RTd��0�h����!
���M,�,�i��E!?RLSYNCFl	�84�!RO�S߸�4��!�
CE��MTCO�M�2�k�)!	��CONS*1�l�u!�WAS�RC|�2�md�!��USB�0�n|�/!STM��'/.�o�Y/��}/p�J/\/�/�/�/�/��I�CE_KL ?%�� (%SVCPRG1�/::$52:???)03b?g?)04�?�?)05�?�?)06�?�?)07OO)0H
TJOE<9ROWK&4 ��O)1,?�O)1T?�O )1|?�O)1�?_)1�? G_)1�?o_)1O�_)1 DO�_)1lO�_Q1�Oo Q1�O7oQ1�O_oQ1_ �oQ15_�oQ1]_�oQ1 �_�oQ1�_'Q1�_O Q1�_wy1%o�/	2)0 ?"0��I1�/�� S�>�w�b�������я ��������=�(�a� L�s���������ߟʟ ��'�9�$�]�H��� l�����ɯ��ۯ��� #��G�2�k�V����� ��ſ���Կ���1���C�g�Rϋ��*_D�EV ���MC:��,����GRP 2��՟�0bx 	�� 
 ,�� ��ߟ���7��[�B� Tߑ�xߵߜ������� ���3�E�,�i�P�� ������z�������� �A�S�:�w�^����� ����������+ O��D�<��� ���'9 ] D��z���� �/h5/G/./k/R/ �/v/�/�/�/�/�/? ??C?*?g?y?`?�? �?�?�?*/�?�?O-O OQO8OuO�OnO�O�O �O�O�O_�O)__M_ __F_�_�?x_�_p_�_ �_oo�_7oo[omo To�oxo�o�o�o�o�o �oE�_i{b �������� �A�S�:�w�^����� ��я�����^+�� O�a�H���l������� ߟƟ����9� �]� D�����z������� �����5�G�.�k�R� ������ſ�����⿀��C�*�<�yϟ�d ���	gϰϛ���`�������+�%�+�<Pߌ����i�� i�y߇�qߧߕ��߹� ����=�"�e���O�=� s�a��������� 3��'��K�9�o�]� �������������� #G5k����� [�W��� C�j�3��� ����/]B/� /u/c/�/�/�/�/�/ �/5/?Y/�/M?;?q? _?�?�?�?�/�?�?�? �?�?OIO7OmO[O�O �?�O�?�O�O�O�O�O _E_3_i_�O�_�OY_ �_�_�_�_�_�_oAo �_ho�_1o�o�o�o�o �o�o�oIooo@o sa�����! �E�9��I�o�]� �������ޏ���� ��5�#�E�k�Y���я ������ן���1� �A�g�����͟W��� ���ӯ	���-�o�T� f��?��������� Ͽ�G�,�k���_�M� o�qσϹϧ����� C���7�%�[�I�k�m� ߵ�����ߥ���� 3�!�W�E�g���ߴ� �ߍ��������/�� S���z���C���?��� ������+m�R�� �s����� E*i�]K� o����/A �5/#/Y/G/}/k/�/ ��/�/�/�/�/�/1? ?U?C?y?�/�?�/i? �?�?�?�?�?-OOQO �?xO�?AO�O�O�O�O �O�O�O)_kOP_�O_ �_q_�_�_�_�_�_1_ W_(og_o[oIoomo �o�o�o	o�o-o�o! �o1WE{i��o ������-� S�A�w�����g�я �������)�O��� v���?�����͟��� ߟ�W�<�N��'�� o�����ɯ���/�� S�ݯG�5�W�Y�k��� ��ſ��+����� C�1�S�U�gϝ�߿�� ύ������	�?�-� Oߥ��Ϝ���u��߽� ������;�}�b�� +��'��������� �U�:�y��m�[��� ���������-�Q� ��E3iW�{� ��)�A /eS����y �u�//=/+/a/ ��/�Q/�/�/�/�/ �/??9?{/`?�/)? �?�?�?�?�?�?�?O S?8Ow?OkOYO�O}O �O�O�OO?O_OO�O C_1_g_U_�_y_�_�O �__�_	o�_o?o-o coQo�o�_�o�_wo�o �o�o;)_�o ��oO����� ��7�y^��'��� �����ُǏ��?�$� 6����W���{��� ��՟���;�ş/�� ?�A�S���w����ԯ ������+��;�=� O���ǯ���u�߿Ϳ ��'��7ύ����� ÿ]Ϸϥ��������� #�e�J߉��}�ߍ� �ߡ�������=�"�a� ��U�C�y�g���� �����9���-��Q� ?�u�c���������� ����)M;q ����a�]� �%I�p�9 �������!/ cH/�/{/i/�/�/ �/�/�/�/;/ ?_/�/ S?A?w?e?�?�?�?? '?�?7?�?+OOOO=O sOaO�O�?�O�?�O�O �O_'__K_9_o_�O �_�O__�_�_�_�_�_ #ooGo�_no�_7o�o �o�o�o�o�o�oao F�oyg��� ��'����� ?�u�c��������� #�����'�)�;�q� _���׏�������ݟ ��#�%�7�m����� ӟ]�ǯ���ٯ��� �u���l���E����� ÿ���տ�M�2�q� ��e���uϛωϿϭ� ��%�
�I���=�+�a� O�qߗ߅߻�����!� ����9�'�]�K�m� ���ߺ��߃������ ��5�#�Y������I� k�E���������1 s�X��!�y�� ���	K0o� cQ�u���� #/G�;/)/_/M/ �/q/�/�/�//�/ ??7?%?[?I??�/ �?�/o?�?k?�?O�? 3O!OWO�?~O�?GO�O �O�O�O�O_�O/_qO V_�O_�_w_�_�_�_ �_�_oI_.om_�_ao Oo�oso�o�o�oo�o �o�o�o']K� o��o���� ��#�Y�G�}���� �m�׏ŏ����� �U���|���E����� ӟ������]���T� ��-���u�����ϯ�� �5��Y��M�߯]� ��q�����˿��1� ��%��I�7�Y��m� �����	ϓ�����!� �E�3�U�{߽Ϣ��� k�����������A� ��h�z�1�S�-���� �������[�@�����$SERV_M�AIL  �����e�OUTPU�Tt���RV� 2�	�  ��� (�O���i�SA�VE��g�TOP1�0 2�� d ��;M_q� ������ %7I[m�� �����/!/3/ E/W/i/{/�/�/�/�/ �/�/�/??/?	��YP��f�FZN_�CFG �	����.��o1G�RP 2�y7�� ,B   A�0~.D;� B�0��  B4.�RB21��HELLr2�	���������7"O1K%RSR1O2ODO}OhO�O�O �O�O�O�O�O_
_C_�._g_R_�_�_�^�/  ��%�_�_P�_�R�\a. �_Lb`ރ��R2. �do�_�6HK 1��; o�o�o �o�o�o�o�o
3. @R{v��������<OMM ���?2��2FTOV�_ENBt����H�OW_REG_U�IR�g�IMIOF�WDL��!��5A���*SYSTE�M*. V8.30�340 ł11/�9/2020 �A ���X�S�NPX_ASG_�T   0 �$ADDRESSo  ��ZE�VAR_NAM	��%$MULTI�PLY��PA�RAM�� � ?$TIME����$�_ID�	�$NUM�D�T�C�IMP[�FRIF�D�VERSION���G�TATU ��$DISK�NFO�D�MODBUS_�ADR[�����POyRC�. �SSR��� x ��N�GLE��g�$D�UMMY7�SG�L�TASK   &����T���<���STMTT0��PSEGT2�BW�D�h��E��SV�CNT_GP�� 8 $PC��ER_V�  _ 	$FB�Pm��SPC��m�ΐVD�X�R[�� �$DATA0ӀS u���1��2��U3��4��5��6��U7��8��9��A��B��C��D��2����F�� y���1Ω1�۩1�1��1�1��1�1)�16�1�C�1P�1]�1j�1Pw�ҁJ���2Ω2۩U2�2��2�2�U2�2)�26�2C�U2P�2]�2j�2w�U3��3��3Ω3۩U3�3��3�3�U3�3)�36�3C�U3P�3]�3j�3w�U4��4��4Ω4۩U4�4��4�4�U4�4)�46�4C�U4P�4]�4j�4w�U5��5��5Ω5۩U5�5��5�5�U5�5)�56�5C�U5P�5]�5j�5w�U6��6��6Ω6۩U6�6��6�6�U6�6)�66�6C�U6P�6]�6j�6w�U7��7��7Ω7۩U7�7��7�7�U7�7)�76�7C�U7P�7]�7j�7w��O͑VPRM_U�PDӑ  9$4q� 
�����ӑؐ$TOR�QUE_CMD �  u�MOa_�SPEEjQ_C�URREo�nAX�I �mS�CAkRT��_Ut�z�͑YSLO�? � ��� ���������_�{�oVALU�OP���$�#(F�ID_�L��K%HIF*IN��$FILE_A�v$�$M�t���SAR0  h�^� E_BLCK����"���(D_CPU�)��)��F#y/�$����_=�R 	� � PWҐO�T��)1LA#�S�R� .3?184RUN_FLGQ5-4U184WITX5v1-4v185�H2�D4�084@�T�BC2��
 �' $O�X0IGu >�0_FTM1D��4]2D�TDCX0AZ���2M���6�1�7T�H��C�DxGRx.0A��ERVE�3�?D�3?D3O��0_A�C@ X ;-$jALEN�3wD��3j@EL_RATmI��$�W_��F#1jAc$2�GMO��!>��C��ERTI�A�o!�Iaj@�KD�E�E��LACEM��CC�CmV�@M�A��F7UW7QTCqV>\_QWTRQ^\ UuZ���Ct��USt��J_��q�M�TF�JH2'���E�QUvA�2�P>�s�a�C@JKfVK�1'a�1'a�`A`J0<d+cJJv3cJJ;cAAL+cPa`3ca`[f4\e5C�PN1�\�`Q[;P��L�@_�E�.�0C�F� `^GRCOU1 ����y�N�0�CC��`REQUI9R*B��EBUZ�fAn�V$T�@2#q�g@v�14 \��ENABL	��$APPRpCL~�
$OPEN`x_CLOSEozSE�y�E
�1.� �u M�0<PPB�t_MGr!�pC��� �x���9P�wBRK�yN�OLD�vh�RTMCO_�3���uJ"��PcdP3cP;cPcP�cP6P��S�>b� ��eB�4� r�B�1����1��PATH ��ӁɃӁ�Hσ0�(p9�W�SCATr�lar�qINiBUC�@���)�C��UM2�Y�@+@�P9�O!EAT���0T�`@T�PAYL�OA�J2L7R'_AN�1��L*0��𛑏����uR_F2�LSHR9DؑLO���(�ٗF��F�ACRL_�!&��"���rBH$ �$H�r^G�FLEXcs�1J�6 PMr�?�?�>OPO�"d�iE :vO�FP٧�O`AP�O�O�LF1� >�R��O�O�O�O_!_��E+_=_O_a_s_�_ �_�_�_Y�vĽW�Sd�f����_�_ o�jT2'W�X�`�eŴ�� e'� �*o<oNo``de me[ee�o�o�o�i�2J�d ��0�o�o� 8ATk�q�PCELٰ}1=�xJ(p�#pJE �CTR�"�f�TNR9�wH�AND_VB��c�0 �� $��Fi2�v	D#SW�!�^�2�v� $$M���yv�q���q �����>��AR ���vQ!5��}A�| �zA�{A�@��{� �zUD�{D�P�G@0���ST�w���y��N�DYW0^p�v!�H� ��k@ϗ�ϗꑎ�g������PX�a�j�`s�|������� Ģ�� ��Ť��x��qASYM��^�p������_�0�.�A�+�-@��K�]�o�����J���K�����˙x�_V�I��	(�s V_�UNIC.$P�בJ eG"uG"�K$�X$ |&
��P�K�,�>��%��T�\��1�0H+0Rr���!v�VrSDI�sO4�1�� �c `�O�I2AO�F�I1l�WW3�o�~0�0ܰ�  o � ��ME���@r2�"YT0P�T���ڀ�1�`�d u���8�1�9T��a� $DUMM�Y1`A$PS_6i�RF+�  ڀ�6�XpFLA�`YP���B�3$GLB_T��5*E�0Vq�`8��j�v1 XMpw֤�ST±#pSB}R��M21_VrT$SV_ER��1O� pC�CCLD@pBeAڰOL2� GL ;EW� 4�`�1W$Y��Z��W�C`ԑ��As02��0�C]U�E ��N�@޵$GIz�}$�A �@�C�@�� L�`V�}$�F�EVNEARʻ�Np�F]Y��TA�NCp��`JOG��A� ��$JOINT
Ѻ`�E�MSET�  "WECU۱�S�'U|��� g��U��?�#pLOC�K_FO���0B�GLVm�GLhT?EST_XMcp�Q'EMP�Pr+bBB��P$U���B2�2#p�CQab���PQarACE�`Sr`_ $KAR�M3TPDRA�@�d�Q�VEC��f�PIU�QaVaHE�PTO�OL2��cV1�REN�`IS3���b6s�Nf�ACH�P(p�a1O��3�429�2�`�ISr  @$R�AIL_BOXEz
��@ROBO"d�?��AHOWWA�RO�Aq�0qROLM�2gu��
txr��/p�Z���O_F��!� �D�a� �_ +�R�`Oˢ!�r*�d�Q�p-2�AOU�R	"XBMeYC���P_$PIP#fN����b/r�ax�Qa�p��CORDED�P��q�� ��OY0 # 7D )@OBu�G� �Pd�S��3(@S��I�wSYSS�ADRH�� �0TCH�S� M,0EN2�A�Q�_T������PV�WVAu1% �� �`�B5PRE�V_RT�$E�DIT�VSHW�R��\F$����A�	 D�0��;���$HEAD�� U����KE�A�0C�PSPDl�JMP�p�L5b�R��44Q&[�t���I,`SH�C��NE�`I��T�ICK2�<M}�۩��HNRA'� @]�����t�_GqP�&v��STY��qLODA,3����m�_( t 
 �GƅS%$�T=\@S>�!$=!2��1EF0rFP�SQU�`x%�B!TERC�0���TS��) Ph@�׹���g��ab�`O�0�3t�IZD4QE�1PRE��1�!����pPU�1�_�DObR��XS�PKN6AXIP��sVaUR�ڳI�Hp�~�d���_�`��ET��QP bl�O�F2P�A�4 s�s`�-2SR��*lѠ��A���� ����#��1�� A�R�c�R�s�RŃ�d� ~Ͱ�dŢ���������C��|�����SC,@ + hƕ@DS��a�0SPLC0~�ATq��2��𐿒�2ADDRE�S�cB�SHIF��H`_2CHH�rz�IK@���TV�I72,��h���� �
+j
�Q��>���- \����O������<�C��򢵲����B<��TXSCR�EEU�.	0k�T�INA�CP��T�np�pQ_��� / T���@����Ag@���^���^����RRO�L wP��f���v�-1UE��0 �� ��@9S�A��RSM�T�UNEX��6F�� S_�Cf�6V�i����6��C�RB��� [2/��UE�1=2��B��!�GMT� L�i!m�w@O�WBB�L_pW�0��2 ��O�O�AL1E��GpTO�3�RIGH&BRD<�D��CKGR�0N�TEX��OJWIDTHs1�u��1AZ�a%�I_�0H�� 3 8�!wP_T��ҭ�0R�@�Rs�w�2$� O�ѭ�4����GG U2 �R brqLUM�u���GERV
���� PaPԒУ5{0�GEKUR&cF���Q)]��LPM��E��C�)�jS�x�x�`w5*u6u7u8Z��@�3�9P��6�a�Q�S��4�USR��D6 <���0U8R��RFOC�aPPRIαmp�!L �TRIP+qm�SUN$0547	Pt��$0��Yq��Hb���� �8�  �G �\�T�p1��ѣ"OS�1�&R���#�a�9�O�C�N�"�$�Ia	UU�:�/�/�U���#OFF!`��;j[�3On0 ٰ�W5�4:�@GUN�w��0B_SUqB�2p@��SRT� ��<��vQ�p �OR�p�5RAU��4T��9���1_���= 9|���OWN� T$SRC���r��D!`CE�MPFI8*�*ё�ESP-��� ���e*B�&�b�!B����> `10WO�8�T�COP&:1$��� _^@�bX�A�q�EWA�C?a��A�@�C�A�b ��VCCH�? ��qC36MFB1����PVC4�Y`��@�x %rT��� XdP^��spC�pRU�DRIV���_�V�uT̐fpD�MY_UBY�ZTV�񕠧�B��X�a�RGP_Sp�+��RL7��BM$��DE�Y��EX����EM�U��X7d[�US�P�po��<1G��P�ACINΑ}�RG MAadwbF3wb3wb���ARE����a�rH6Twb�pA R�@G�P�Pr�a6UR� �pBC d�_���2	�B�N�RECcSWo`_IApa�8c�O!���A��1s�E�U`B�� �q�8SHKG�C��Iz���.p��zsEA���w�@� 1u�5UMRCV��D U�FOS�M� Cs��	�rX3�c�rREF ���v�v�q p7��p  �z��z��{;��v�p_@@�zq��{��S��/g�S�6�8R��E �$�=�ߠ) �UӠOU��b�ZSO @�e2�2�a$��R� �ΐB��t2Ѻ�Kq�SULs��C�@CO:�� D)`�NT�CZ�R@Y��e�!e�$�L�S����S�����!�|JTǤFt +���ǱT� ��CACH+�LO����*`�����@ܣC_LIM-I��FR%�Tj�'�N��$HO� 6B�OCOMMpSB�O0 �]�Ԉ�I؄h@VPx�bP��_SZ3n�2��6����12����[`��&����AaMP��FAI&�Gvt���AD��BMRE�ׄ9�_SIZ�P�H�`��FASYN�BUF�FVRTD�k�w�I�aOL��D�_@3��W3P�E�TUc�QNp[�EwCCU�hVEM�`x��۲&�VIRC���VTP�pO��J��s�A�w�_DELA��cP�Ʃŕ��G��@9pCKLAS��3	ő_�F�ƀH$p"�S;��N��P/LEXEEI��B�/��3cFLK I  `]�^A��M���dws�Yr/�^@�bJ# ��ʱ��#�#RS ORD@!�4Q> 3 ނ�)�K��T\"����WwCb2V��g%L`�Qۑ6D4��\*b3UR3cp_R'�d� ��,a]��ծc�_od@&�{g��`B*�T�N'�SCO��*�C�  ad�"_f�"0�">�" K�"Y�J_\_nZ���� E\ AM�P�0� PSMf%M�p"%HADJT�/e��Bڒ� Np"q׬!�LIN]3q��XV�Rh$O\���T_O�VR� �ZAB�C�5P�bw�$��
���ZIPg%Qp"D/BGLV�CL�R �}�ZMPCF�5GR  r ���$��.�QLNK�2
��-`�|�S �|q����CWMCMi`C�CC�A�CtP_�  '$J:4D��@ QJ�V�4$0�t�O�UXW� ��UXE>a��E�[����	��u���T ����r�Y:K�D"0 U�"�֝^IGHbcq�?�( �K��V� � vG��$B�$��@1e�B�҉�&GR�V%�F� ���OVC�5�A7�w@�`�J�
VBI���D�_TRACEB�V;1}�SPHER�P W , �3I>[�$SIM�A�!82Re!�� �e!V&��qe!�m/!��%����/Kpb/t#_sUN�@_+p&�LCд�% �%�V M��ALIAS ?e���%1~�! ( he�! :?L?^?p?�?�66?�? �?�?�?�?	OO-O?O QO�?uO�O�O�O�OhO �O�O__)_�OM___ q_�_._�_�_�_�_�_ �_o%o7oIo[ooo �o�o�o�oro�o�o !3�oWi{�8 �������/� A�S�e���������� я|�����+�֏<� a�s�����B���͟ߟ ����'�9�K�]�o� �������ɯۯ���� �#�5��Y�k�}��� ��L�ſ׿���ϸ� 1�C�U�g�y�$ϝϯ� ����~���	��-�?� ��c�u߇ߙ߫�V��� ��������;�M�_� q��.�������� ��%�7�I���m�� ������`������� !��EWi{&� �����/ AS�w���� j��//+/�O/ a/s/�/0/�/�/�/�/ �/�/?'?9?K?]?3��$SMON_D�EFPRO �����1� *SYS�TEM*p:REC�ALL ?}�9� ( �}2xc�opy fr:\�*.* virt�:\tmpbac�k�1=>172.�8.9.225:?14224 �2�?XO!O2M}3�5a�?��?�4�?�O�O�OB@7��4s:orderfil.datTL`fO|O__1_}.�2mdb:QO�Ox@�O �_�_�_>D�?XO�?{_ oo0oCO�_�_yO�o �o�o�O�O\_w_ ,?_Q_�o�o��� �_Pobo�_��(�;o�Mo�qo������9�
�xyzrate 11 Q�c�u����*�=�Ƈ�8644Ё������������Q�c�u���*�=�|F��t0836 � ���������o�oYZ� ���!�4F�Y����������=�Ưبem=p`}680 z����/�B�+ƶ*.d ڿ��ϕϧ�:�L��m�d�v���+�>�:��th:\supp�ortP�P�=>4�79854592?:64327�ϐ���5��qՃoutp�ut\untitled8.pcJ�?: overm�� �"������9���������;�tpd_isc 0�� a��s���(�;�tp?conn 0Л�� ��2�������ȆQ�c��u�*��O�7252 ������� ��Qas(;��M���2��6�9�F���1��3519�2832]�268�8�/"/����2����/�/�/;���35�pd/v/??+?>���'�/�/�?�?�? <N�]?o? OO$O7? I?�?�?2O�O�O5O�3 �/_OqO__&_9OKO �O�O�_�_�_�?�?[_ m_�_o"o5/G/��]69752o�o�o��ǿٯ�_ ~o!4� F��o�(�o���;���$SNPX_A{SG`����q�� P �0 '%R[1]@1.1��y?�;�%�(�� L�/�A���e������� ܏��я����H�+� l�O�a�������؟�� ��ߟ�2��<�h�K� ��o���¯��̯��ۯ ����R�5�\���k� �������ſ���� <��1�r�U�|Ϩϋ� �ϯ�������8�� \�?�Qߒ�uߜ��߫� ������"��,�X�;� |�_�q�������� ����B�%�L�x�[� ������������� ,!bEl�{ ������( L/A�e��� ���/�/H/+/ l/O/a/�/�/�/�/�/ �/�/�/2??<?h?K? �?o?�?�?�?�?�?�? O�?ORO5O\O�OkO �O�O�O�O�O�O_�O <__1_r_U_|_�_�_ �_�_�_o�_o8oo \o?oQo�ouo�o�o�d��tPARAM ��u�q ��	��jP;tAp��h#t��pOFT�_KB_CFG � s�u�sOPI�N_SIM  �{vu��p�p�RVQSTP_DSB^~r��x�`�SR ay �� & SOCgKET�"��v�TOP_ON_ERR  -�Kx?�_PTN �fr��A;�RIN�G_PRMI� ��`VCNT_GP� 2au&q�(px 	�̏p���ޏ���wVD��RP 1�i'p�y� R�d�v���������П �����*�<�N�`� ����������̯ޯ� ��&�M�J�\�n��� ������ȿڿ��� "�4�F�X�j�|ώϠ� ������������0� B�T�f�xߟߜ߮��� ��������,�>�e� b�t��������� ���+�(�:�L�^�p� ��������������  $6HZl~� ������  2DV}z��� ����
//C/@/ R/d/v/�/�/�/�/�/ �/	???*?<?N?`? r?�?�?�?�?�?�?�?�OO&O0�PRG_�COUN�At�8r�NuRBENB��ME�MwCAt�O_UPD� 1�{T  
;Or�O�O�O__ (_:_c_^_p_�_�_�_ �_�_�_�_ oo;o6o HoZo�o~o�o�o�o�o �o�o 2[V hz������ �
�3�.�@�R�{�v� ����Ï��Џ��� �*�S�N�`�r����� �����ޟ��+�&� 8�J�s�n��������� ȯگ����"�K�F� X�j���������ۿֿ ���#��0�B�k�f��x�DL_INFO {1�E�@��	 ����������@L�g@�D��?��{��	
� �	̀���@������%^��ຏA�f��o߁�� D��D��q}D�Q�6���p´�ߞ�O@Y?SDEBUG\@�@���d�I��SP_�PASS\EB?~��LOG �ƕ�C���ؘ� � ��A��UD�1:\���_M�PC�E���A�H�� �Am�SAV �m�4�L���S�SVd�TE�M_TIME 1u	��@ 0���R��P��_��$T1SVGUNS�@�]E'�E�r�AS�K_OPTION�\@�E�A�A��_D�I��xO��BC2_?GRP 2
�I=�|��Ѡ  C��f�BCCFG ����� l�]`]`ߕ��� ����7"[ FX�|���� ��/3//W/B/{/@f/�/�/�/�/���, �/�/"?4?�/?j?U? �?y?�?���?���0�?  O�?$OOHO6OlOZO |O~O�O�O�O�O�O_ �O2_ _B_h_V_�_z_ �_�_�_�_�_�_�_.o h� BoToro�o�oo �o�o�o�o�o&8 \J�n��� ����"��F�4� j�X�z�����ď��� ֏�����0�f�T� ��@o����ҟ���t� ��*�P�>�t����� f������ί��� �(�^�L���p����� ʿ��ڿ ��$��H� 6�l�Z�|�~ϐ��ϴ� �Ϡ���2�D�V��� z�hߊ߰ߞ������� ���
�@�.�d�R�t� v����������� *��:�`�N���r��� ������������& J �bt���4 ����4FX &|j����� ��//B/0/f/T/ �/x/�/�/�/�/�/? �/,??<?>?P?�?t? �?`�?�?�?OO�? :O(OJOpO^O�O�O�O �O�O�O _�O$__4_ 6_H_~_l_�_�_�_�_ �_�_�_ ooDo2oho Vo�ozo�o�o�o�o�o 
�?"4Rdv�o �������� �<�*�`�N���r��� ����ޏ̏���&�� J�8�Z���n�����ȟ ���ڟ�����F�4� j� ������į֯T� ���
�0��T�>�r���$TBCSG_�GRP 2>���  ��r� 
 ?�  ������ӿ����῀�-��Q�c�v�}�~��d0 ����?r�	 HC��`�r���b�C�  �B����Ȣ�>�ff�źƞ�����)��϶�\��H �hݳBLcφ�B$д h�j߈ߎ߲߰�����	���@�@��AƷ�f� y�D�V��������	��?333���2�	V3.00~��	m2ia�	*T�L�q�c�"�.���r������ ��l���   ��B������u�J2}���5����CFG >�e�� ��
�D9��o�o� �
G������ �5 YDV�z ������/1/ /U/@/y/d/�/�/�/ �/�/�/�/????Q? ����\?n?�?*?�?�? �?�?�?O�?1OOUO gOyO�OFO�O�O�O�O �O	_r�^�._:�>_@_ R_�_v_�_�_�_�_�_ �_o*ooNo<oro`o �o�o�o�o�o�o�o 8&\Jl�� ��������� 6�X�F�|�j�����ď ��ԏ����܏.�0� B�x�f�������ҟ�� �����*�,�>�t� b����������ί� ��:�(�^�L���p� ������ܿʿ ��$� �H�6�X�~�(��Ϩ� ��d����������D� 2�h�Vߌߞ߰��߀� ����
����@�R�d� �t��������� �����*�`�N��� r������������� &J8n\~� �����"�� :L
�|�� �����0/B/T/ /d/�/x/�/�/�/�/ �/?�/,??P?>?`? �?t?�?�?�?�?�?�? OOOLO:OpO^O�O �O�O�O�O�O�O_ _ 6_$_Z_H_j_l_~_�_ .�_�_�_�_ oo0o VoDozoho�o�o�o�o �o�o�o
@.P v��Tf��� ���<�*�L�r�`� ��������ޏ̏��� �8�&�\�J���n��� ����ڟȟ���"�� F�X�op���o>�į ���֯����B�0� f�x���H�Z������ ҿ��,�>���b�P� r�tφϼϪ������ ��(��8�^�L߂�p� �ߔ��߸�������$� �H�6�l�Z��~�� �����d����&��� ��D�V���z������� ����
.��R@ bdv����� �*N<^` r������/ /$/J/8/n/\/�/�/ �/�/�/�/�/?�/4? "?X?F?|?�?8��?�? �?t?�?�?OO.O0O BOxOfO�O�O�O�O�O��O�O__>_(^  9dPhS hV|_�hR�$TBJOP_GRP 20U��  �?�hV	�R�S��\�8P���p��Q�U � � � � y��RhS @dP��R	 �C� >ff  C�W�Q�4b��<f9o >��ff\a<a=�ZwC�`���b�&`H&`.g�o�g�nѴW4e\e`b�o �?a�d=�7LC��noBȂo#&`�p`9u�o�c�33\u�X2h�P<��C�\vc@333@�33|b}`�BL��wHqDa�l����u�Jh�p<X���B$�d��?_���C*p���C���Z`y�x��k<G ��q`?]`�C4.�ϏR�d��da�G����{<gș��]p@&b`yap�c�z{4ep�V� ���������ʟ��� (�� �N��Z����@������ޯ��d�hV�0�4e	V3.�00�Sm2ia�T*Z��TcQh�s�� E�'E��i�FV#F�"wqF>��F�Z� Fv�RF��~MF���F����F��=F����F�ъF���3F���F��{G
G�dG�G�#
��D���E'
EMK�E���E�ɑ�E�ۘE���E���F���F��F���F(��F5���FB��FO���F\��Fi���Fv��F��v�F�u�<#�
/<t���@Ť�Ar_X�j�M�hTn��@�U�S��SESTP�ARSA�\X�P�SH�R��ABLE 1%�[��hS�ȃ�Q �0cɞ����ȨgWoQ��	��
�������hQ����8��C���RDI�ϬQ��� �2�D�Vվ�O����������*���S�ߪS ������ �!�3�E�W�i�{��� ������������ /A�]�����̂	k� }���M�_�q߃ߕ������hNUM  �0U�Q�P�pP B�C���_CFGG P�a@�P�IMEBF_TT�����S���VER�AÔ��R 1=�[ 8e�hR�cP! 3P�   � //$/6/H/Z/l/ ~/�/�/�/�/�/�/�/ ? ?2?{?V?h?�?�? �?�?�?�?�>��?O�:0OBOTO.OxO�O dO�O�O�O�O�O�O_ ,__P_b_�8�_�_ �_~_�_�_�_�_����_K�@���M�I_CHAN� �� mcDBGLV�逡���p`ET�HERAD ?*���`�n��?o��o�o��p`ROUT6�!p
!"t@~|SNMASK�h|��a255.~u�F�|��F���OOLOFS_DI���GT �iORQC?TRL p	��	n��T�B�T�f� x���������ҏ��� ��,�>�P�b�r��𕟄�����PE_D�ETAI�h�zPG�L_CONFIG� Qa���/cell/$C�ID$/grp1���3�E�W�i�{�1� 	����ʯܯ� ��� $�6�H�Z�l�~���� ��ƿؿ�������2� D�V�h�zό�ϰ��� ������
ߙ�.�@�R� d�v߈��)߾���������}��N�`� r��������������)�;�M�_� �߃�����������l� %7I[m�� ������z !3EWi��� ������/// A/S/e/w//�/�/�/ �/�/�/�/?+?=?O? a?s?�??�?�?�?�? �?O�?'O9OKO]OoO �OO�O�O�O�O�O�O�_��User View !��}}1234567890B_T_f_x_��_�_�T-`��_��(Y25Y�Ooo*o<o No`o�_�_/R3�_�o �o�o�o�ogo)�^4�obt������^5Q�(�:�@L�^�p�����^6� ʏ܏� ��$���E��^7��~�������Ɵ؟7����^8m�2�D��V�h�z���럭��� �lCamera3Z)����(�:�L�*�E�v��� ��@_��ƿؿ�����  ̦�Y�^�p� �ϔϦϸ�_����� � K�$�6�H�Z�l�~ߥ��̦�i������� � �$���H�Z�l�ߐ� ���������ߣ�Py ��6�H�Z�l�~���7� ������#��� 2 DV���*����� ������"4F �j|����k ͥ��Y/ /2/D/V/ h/�/�/�/��/�/ �/
??.?���l��/ z?�?�?�?�?�?{/�? 
OOg?@OROdOvO�O �OA?�� �1O�O�O
_ _._@_�?d_v_�_�O �_�_�_�_�_o�O�G9�_GoYoko}o�o�o H_�o�o�o�_�o1�CUgy�	Υ0 �o�������o 2�D�V��oz������� ԏ{�Ӡիx�-� ?�Q�c�u���.����� ϟ����)�;�M� �ΥA�䟙�����ϯ �󯚟�)�;���_� q���������`��u�� P���)�;�M�_�� �ϕϧ��������� �%�̿޵���q߃� �ߧ߹���r����� ^�7�I�[�m���8� ޵�(�������%� 7���[�m������� ����������޵��� I[m��J�� ��6!3EW<i  	� �����//(/x:/L/^+   n v�/�/�/�/�/�/ ? ?$?6?H?Z?l?~?�? �?�?�?�?�?�?O O 2ODOVOhOzO�O�O�O �O�O�O�O
__._@_ R_d_v_�_�_�_�_�_�b,  
 (  ��( 	  �_oo:o(o^oLo�o po�o�o�o�o�o �ot$�Z~* ̸ i{� ���� ��X5�G�Y�� }�������ŏ׏��� ��f�C�U�g�y��� �����ӟ�,�	�� -�?�Q�c��������� �������)�;� ��_�q���ʯ����˿ ݿ��H�%�7�Iϐ� m�ϑϣϵ���� � ���!�h�E�W�i�{� �ߟ���������.�� �/�A�S�e�߉�� ������������+� r��a�s�������� ������J�'9K ��o����� ��X5GYk }������0 //1/C/U/g/��/ �/�/��/�/�/	?? -?t/Q?c?u?�/�?�?��?�?�?�?:?p@ AB"O4OFOCG� `��)frh:�\tpgl\ro�bots\m20�ia\arc_m�ate_1�@c.xmlO�O�O�O�O��O__(_:_L_XX��X_}_�_�_�_�_�_ �_�_oo1oCoZ_To yo�o�o�o�o�o�o�o 	-?VoPu� �������� )�;�RL�q������� ��ˏݏ���%�7� N�H�m��������ǟ ٟ����!�3�J�D� i�{�������ïկ� ����/�F�@�e�w� ��������ѿ������+�=�_H�1 �Oj@88�?�=�|�=�xϚϜ� ���������0��<� f�P�rߜ߆ߨ��߼�����&��$TPG�L_OUTPUT� "H1H1 `�H�]�o�� ������������� #�5�G�Y�k�}����������������H�`����2345678901 2DVh z�>2���� ��9K]o�}����� ���1/C/U/g/y/ �/#/�/�/�/�/�/	? �/???Q?c?u?�?? 1?�?�?�?�?OO�? %OMO_OqO�O�O-O�O �O�O�O__�O�OI_ [_m__�_�_;_�_�_ �_�_o!o�_/oWoio {o�o�o7oIo�o�o�o /�o=ew� ��E�����+�� �}[�a�s���������̍@b�����h� ( 	  7�%�[�I��m��� ������ǟ���!�� E�3�i�W�y�����ï ���կ�����/�e�S����^�w� ��ѽ�����)�;� ��d�v�ϚϬϊ� ����L���ߺ�(�N� ,�>߄ߖ� ߺ���n� �����&�8��D�n� �^��������V� �"���F�X�6�|��� ��z�����x����� 0B��fx�� ���N`,� Pb@���� p�/�/:/�� p/�/$/�/�/�/�/�/ X/�/$?�/4?Z?8?J? �?�??�?�?z?�?O �?2ODO�?POzOOjO �O�O�O�O�ObO_._ �OR_d_B_�_�__�_ �_�_�_oo�_<oNo�Tb�$TPOFF_LIM ���p�����qibNw_SVm`  ӄ�jP_MON �#���d�p��p2ӅiaSTRT?CHK $��f�^��bVTCOM�PAT�hq�fVW�VAR %�m\Ax�d �o Y��p�bia_DEFPROG 3v�b%SOCKE�p��m_DISP�LAYt`�n�rIN�ST_MSK  ��| �zINU�SER�tLCK���{QUICKM�ENA��tSCRE�`���rtpsc�t�{���b���_��STziR�ACE_CFG �&�iAtx`	�bt
?�܈HNL 2'�i}� �H{ nr4�F�X�j�|���𠟲�ĚޅITEM� 2( � �%�$1234567�890��  =�<�7�I�Q�  !W�_�kp���bs �ů)����_���� ��^���y�ݯ����5� %�7�I�c�m�翑�=� c�u�ٿ�����!ϛ� E����)ߍ�5߱��� ��Yߧ������A��� e�w�@��[���� �ߧ��k���O��s� �E�W���c������ }�'�����o�/�� ����;S����# �GY"}=�a s����1� U/'/����� �_/	/�/�/�/Q/? u/�/�/?�/i?�?�? ?�?)?;?M?�?O�? COUO�?aO�?�?�OO �O7O�O	_mO_�O�O l_�O�_�O�_�_�_3_ �_W_i_{_�_�_Koqo �o�_�ooo/o�o�o eo%7�oC�o�o� �o���O�s(�N�ڄS�)�S���  ϒS�q �����y
 ���ݏď���UD1�:\���e�R_�GRP 1*��� 	 @�p Y�k�U���y�����ӟ�������͑�2�x�V�A�?�  q� ��m�����ǯ���ٯ �����E�3�i�W���`{��������	!�����c�SCB 2+o� \�Y�k� }Ϗϡϳ�������Y��V_CONFIG ,o�󁧏�M����OUTPUT �-o�>��� Yߝ߯���������	� �-�?�Q�c�u�;ъ� �����������	�� -�?�Q�c�u������ ��������); M_q������ ��%7I[ m������ �/!/3/E/W/i/{/ ��/�/�/�/�/�/? ?/?A?S?e?w?�/�? �?�?�?�?�?OO+O =OOOaOsO�O�?�O�O �O�O�O__'_9_K_ ]_o_�_�O�_�_�_�_ �_�_o#o5oGoYoko }o�_�o�o�o�o�o�o 1CUgy� '�9Ո������ #�5�G�Y�k�}����� �oŏ׏�����1� C�U�g�y��������� ӟ���	��-�?�Q� c�u���������ϯ� ���)�;�M�_�q� ��������˿ݿ�� �%�7�I�[�m�ϑ� �ϴ����������!� 3�E�W�i�{ߍߟ߱� ����������/�A� S�e�w������� ������+�=�O�a� s��������������� '9K]o� �������� #5GYk}��|��x���� ���/�3/E/W/ i/{/�/�/�/�/�/�/ �/?�/?A?S?e?w? �?�?�?�?�?�?�?O O*?=OOOaOsO�O�O �O�O�O�O�O__&O 9_K_]_o_�_�_�_�_ �_�_�_�_o"_5oGo Yoko}o�o�o�o�o�o �o�o0oCUg y������� 	��,?�Q�c�u��� ������Ϗ���� (�;�M�_�q������� ��˟ݟ���%�6� I�[�m��������ǯ ٯ����!�2�E�W� i�{�������ÿտ������,��$TX�_SCREEN �1.����}ipnl�/`�gen.htm,�ϑϣϵ���$ �Panel �setup��}������0�B�T�f� ���ϝ߯��������� n���?�Q�c�u�� ���"��������� )�������q������� ����B���f�%7 I[m������� ���t��EW i{���:���////A/�/�U�ALRM_MSG� ?L��Y�  Z//��/�/�/�/�/�/ ??$?B?H?y?l?�?��?�?u%SEV  ��-�6s"EC�FG 0L��V�  /�@� � A#A   B�/�
 �?6�L�VO hOzO�O�O�O�O�O�O��O
_W�1GRP �21	K 0/�	� @Ob_u I_B�BL_NOTE �2	JT�G�l6�Q�8�@~uRDEFPRO =%�+ (%�?�_ 8��_o�_'ooKo6o ooZo�o�o�o�o�o�o�k\INUSER � �]P_�oI_M�ENHIST 1�3	I  ( ��P��(/SO�FTPART/G�ENLINK?c�urrent=m�enupage,153,17������'q�~71@�+�=�O�a��q+�ރuedit�rSOCKET���ŏ׏ f��o��1�C�U�g� ����������ӟ�t� 	��-�?�Q�c��� ������ϯ�󯂯� )�;�M�_�q�<x�Rlq �����Ϳ߿��� '�9�K�]�oρ�ϥ� ���������ώϠ�5� G�Y�k�}ߏ�߳��� ��������1�C�U� g�y���,������� ��	����?�Q�c�u� �������������� ),�M_q�� �6���% 7�[m��� D���/!/3/� W/i/{/�/�/�/�/R/ �/�/??/?A?�/e? w?�?�?�?�?�����? OO+O=OOOR?sO�O �O�O�O�O\O�O__ '_9_K_]_�O�_�_�_ �_�_�_j_�_o#o5o GoYo�_}o�o�o�o�o �o�oxo1CU g�o������ �?�?�-�?�Q�c�u� x������Ϗ�󏂏 ��)�;�M�_�q���� ����˟ݟ����%� 7�I�[�m��� ��� ǯٯ������3�E� W�i�{������ÿտ��������$U�I_PANEDA�TA 15����A�  �	�}/fr�h/cgtp/w�holedev.stm�{ύϟϱ�>��)prii�����}���"�4�F�X�j� )lߐ�wߴߛ� ���������2�D�+�h�O�������  � O����� #�5�G�Y���}��ϡ� ����������b�1 U<y�r�� ���	�-?&c�� D��CÞ�� �����P!/�� E/W/i/{/�/�//�/ �/�/�/�/?/??S? :?w?^?�?�?�?�?�? �?Oz�=OOOaOsO �O�O�?�O./�O�O_ _'_9_K_�Oo_V_�_ z_�_�_�_�_�_o#o 
oGo.oko}odo�oO &O�o�o�o1�o Ug�O����� �L	��-�?�&�c� J������������� ڏ���;��o�o~�� ������˟ݟ0��t %�7�I�[�m��柣� ����ٯ�������3� �W�>�{���t����� տ�Z�l��/�A�S� e�w�ʿ��������� ����+ߒ�O�6�s� Zߗߩߐ��ߴ���� ��'��K�]�D���� Ϸ����������d� 5�G���k�}������� ��,�����C *gy`�����������}��,ew����) S�W��/"/4/F/ X/j/��/u/�/�/�/ �/�/?�/0?B?)?f? M?�?�?�?�?Q������$UI_POSTYPE  ���� 	 ��?#O�2QUICKMEN  K�O&O�0REST�ORE 16���  �	�?X��O�C�OX�m�O�O__'_9_�O ]_o_�_�_�_H_�_�_ �_�_o�Oo0oBo�_ }o�o�o�o�oho�o�o 1C�ogy� ��Zo���R� -�?�Q�c�������� ��Ϗr����)�;� ���Z�l�ޏ����˟ ݟ����%�7�I�[� m��������ǯٯ�� ���
�|�E�W�i�{� ��0���ÿտ���π��/�A�S�e�w�1GS�CREA@?FM�u1sc�@�u2��3��4��5*��6��7��8���2�USER���ϫ�TL����ks���4�U5�6�7�8���0NDO_CFG� 7K<;�0P�DATE �����ޝ4B���_INFO 1e8����RA0%}� ��Q��������'�
� K�]�@��d������������*L��OFFSET ;FM�Ë@ �b�t��� ������������N� UL^����@���&VO(
�L*�UFRAME�  �d֑�R�TOL_ABRT8p�ӈENB��?GRP 1<�IRACz  A�� ����	//-/?&!I/[/�@@U�i�~�MSK  ���ӢNm%��%x��/�_EVN�b�$c�
6U�2=I�9hi�UE�V�!td:\�event_usger\�/T0C7Y?d)�F�<L1SPR1�W7spotwe{ld�=!C6�?�?�?�@�$!�/h?&O [OGl�OJO8O�O�O nO�O�O�O_�O�O�O e__�_4_F_|_�_�_ �_�_�_�_=o,oaoo o�oBo�o�oxo�o�o'�o�j)6WRKg 2>@�88"�� y���� 
��.�@��d�v�Q� ������Џ⏽�����<�N�)�_�������$VCCMU�?l\ݨ�MR�2E8;�<�"�	j����~XC56 �*����h� ��5�i�A@7 p:? ȗ� ;[�e�Ȇ���ů�����^�9%A���ٯ*�� B���E��I�ѯj��� ��]�����ֿ����� ��0χ��f�Q�cϜ��O����ϥ�ISIO�NTMOU? ���ů�FU���U�(� �FR:\��\u�A��?  �� �MC*�LOG7� �  UD1*�E�X[�E!' B@ ����o�r���o������d ��  =	 1-� n6  -����Ҭ6,�ր�1�O=���:���n�}P�TRAIN�� ��1�E!�Ad��͓G8; (��:�� S�����������-�� 1�?�Q�c�u��������T���_��RE��Hx�����LEXE���I8;�1-e��V�MPHASE  ����A���RT�D_FILTERw 2J8; ��R������� 1C#��t� ������//���SHIFT�"1K8=<���/p/3��O/u/�/�/�/�/ �/�/?�/?)?b?9?�K?�?o?�?�?�?	�LIVE/SNA�P�3vsfli�v4�?��� �SETU�0BmenuOO�?}O�OfBl/%L���	|H�{O�O��?�J� ��@-�AdB8��B���K�M�QR�S�����	'-_MEh�0�ļ�/!MO�M �zWqWAITDINEND�����TOK  �噰\���_S�_�YT�IM����
lG �_,m�_Ok�_/j�_/j<o�XRELEK_g྘�Q��֗Q_AC�T�0^h(q�X_3� N��)r%�O_���rRDIS�0�n_�$XVR�BO ��$ZABC͒1�P�� ,����2\g7ZIP�CQ�����/�A�S��zMPCF_G 1R�J��0��w��a�MPb�sS���<������8�����3̟�?��  �����w�ȿ������D��D�q_}D�Q���?�����:��hK�=�&7��);��=>�T�d��(�:�;B�T�f� v�e�Ο����A�2�?6��p´$�6� >Ȇ�n�h�z�����ȫ��pt��T|��w�Y�LINDqU|��  �e� ,(  *)�:���&�c�J���n� ���Ͽ� #��s�(��!�^ϡ� �ϔϦ����e�K� � ��$��y�Z�l��{��s2V�+q đ� �������������h��D��ז^�A����SPHERE 2W	�̾Ϛ�ߓ��� ����<�O�*�<���`� �����}�������� I�[�8��\CU��������pZZ�f ��f