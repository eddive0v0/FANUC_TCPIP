��  I��A��*SYST�EM*��V8.3�0340 11�/9/2020 A   ����SBR_T �  | 	$S�VMTR_ID � $ROBO�T9$GRP�_NUM<AXIaSQ6K 6NFF�3 _PARAM�F	$�  �,$MD SPD�_LIT  &2�*  � �����$$CLA�SS  ���������� V�ERSION��  ��~�IRTUAL���'  1 �� T���A�RC Mate �120iC���  �aiS12�/4000 80�A��
H1 D�SP1-S1��	P01.05W,  	� v���  ��# :�����������{  ���r9 � �9����� HH��  �����
/m����  D�4�Z %u%����� ����� 1��2M��?�X���B=��d�����&���<
= z ���� J�����������; � �����T���N��.���Y	�?  � !�� �� :?8���?'by�c/�/0�/�/?��?;?�!R?d?v?�?��2�/1��>���x���r��2*->�0�����o��>�?�?�I�<N`r2|�2�� ��� } J  	����^�,������A �'/ӹ/�A#�"p�< 2�"t���=��	���7_��
��D<)�J �� ���� ErV$��?p$��z(w>��q"��P�(�/�/���/�_�_�_ �_ ?�_D?oo1oCo�0�"��@�����
P,$b�b3dH�@~������:�3�uFo�o�T\�?N@8NJw3|3<ONI
[K_&������wB
=� �D���S�J8H�B ,P����.��+{ ]'H�H�&�����1�/����>��� �� �23
���KvB� ���
P�@X"��op# ���Z 2|%j���  ��l�&WBVR� d~^Sc A�jS{:rY:q� K�]�o����_����� ҏ�����,�>����ɬoNbV@/6!A4�k4|�b�o���P���ϓp�`�M������{���99�� ���"@D@�r�[ ��X"�� �'��sBC�U�~��� 	�����,V$y���  ��� ��s;@2���q"�� �D��%����p(�����'jT�rYT� ����'�9���]��� ��������ɿۿ���rZ��d�N��	R��x5|�b��.Ԛ�������X � ��/X"�� ��!-�?��������*�p$qP�r��1��zR��Q ��&�į֯诱��� ����B��f�/�A�S��e�w��������N@�r6|6�d�v�О����YҨ�� ��2�X"��Q���������-�����t ���!����qTa
��#�&�|ߎߠ� i{������� �/ASew�������xTa��Ng�	�LA���/ / 2/D/V/h/z/�/�/�/ �/�/�/�/
??.?@?P<�P?t?�?�?�?�? �?�?�?OO(O0C� �FO����O�O�O �O�O__*_<_N_`_ r_�_�_�_�_�_�_�_ o^?&o8oJo\ono�o �o�o�o�o�o6OhOZO #~O�OXj|�� �������0� B�T�f�x�������
o �������,�>�P� b�t������o����* <N�(�:�L�^�p� ��������ʯܯ� � �$�6�H�Z�l�ȏ�� ����ƿؿ���� � 2�D�V�ҟğn���� �������
��.�@� R�d�v߈ߚ߬߾��� ������*N�`� r����������� �^ϐς�K��ϸπ� �������������� "4FXj|�� ���2��0 BTfx���� ���R�d�v�>/P/ b/t/�/�/�/�/�/�/ �/??(?:?L?^?p? �?�?��?�?�?�? O O$O6OHOZOlO~O� ��O/"/4/�O_ _ 2_D_V_h_z_�_�_�_ �_�_�_�_
oo.o@o Ro�?vo�o�o�o�o�o �o�o*�O�O�O s�O�O����� ��&�8�J�\�n��� ������ȏڏ���Zo �4�F�X�j�|����� ��ğ֟�D� �z ��f�x��������� ү�����,�>�P� b�t����������� ���(�:�L�^�p� �ϔϦ�"����8�J� \�$�6�H�Z�l�~ߐ� �ߴ���������� � 2�D�V�h�z�ֿ��� ��������
��.�@� R������ϛ������ ����*<N` r������� &��8\n� �������/ l�5/(/�������/�/ �/�/�/�/�/??0? B?T?f?x?�?�?�?�? �?�?@OO,O>OPO bOtO�O�O�O�O�OJ/ </�O`/r/�/L_^_p_ �_�_�_�_�_�_�_ o o$o6oHoZolo~o�o �o�?�o�o�o�o  2DVhz�O_�O �_0_�
��.�@� R�d�v���������Џ ����*�<�N��o `���������̟ޟ� ��&�8��]�P�� ����ȯگ���� "�4�F�X�j�|����� ��Ŀֿ����h�0� B�T�f�xϊϜϮ��� ������r�d�߈��� ��t߆ߘߪ߼����� ����(�:�L�^�p� �������&��� � �$�6�H�Z�l�~��� ����0�"���F�X�  2DVhz��� ����
.@ Rdv����� ��//*/</N/`/ ���/x/���/�/ ??&?8?J?\?n?�? �?�?�?�?�?�?�?O "O4O�XOjO|O�O�O �O�O�O�O�O__�/ �/6_�/�/�/�_�_�_ �_�_�_oo,o>oPo boto�o�o�o�o�o�o �oNO(:L^p �����&_X_J_ �n_�_H�Z�l�~��� ����Ə؏���� � 2�D�V�h�z������o ��ԟ���
��.�@� R�d�v��������� ,�>���*�<�N�`� r���������̿޿� ��&�8�J�\ϸ��� �Ϥ϶���������� "�4�F�¯��^�د� ������������0� B�T�f�x������ ��������v�>�P� b�t������������� ��N߀�r�;�ߨ�p �������  $6HZl~� ���"���/ / 2/D/V/h/z/�/�/�/ �/�/BTf.?@? R?d?v?�?�?�?�?�? �?�?OO*O<ONO`O rO�O��O�O�O�O�O __&_8_J_\_n_�/ �/�_ ??$?�_�_o "o4oFoXojo|o�o�o �o�o�o�o�o0 B�Ofx���� �����v_�_�_ c��_�_������Ώ�� ���(�:�L�^�p� ��������ʟܟ�J  �$�6�H�Z�l�~��� ����Ưد4����j� |���V�h�z������� ¿Կ���
��.�@� R�d�vψϚϬ���� ������*�<�N�`� r߄ߖ�����(�:� L��&�8�J�\�n�� ������������� "�4�F�X�j��ώ��� ����������0 B�����ߋ����� ���,>P bt������ �//r�(/L/^/p/ �/�/�/�/�/�/�/ ? \%??���~?�? �?�?�?�?�?�?O O 2ODOVOhOzO�O�O�O �O�O0/�O
__._@_ R_d_v_�_�_�_�_:? ,?�_P?b?t?<oNo`o ro�o�o�o�o�o�o�o &8J\n� ��O������ "�4�F�X�j��_�_�_ ��o o�����0� B�T�f�x��������� ҟ�����,�>�� P�t���������ί� ���(���M�@��� ̏ޏ����ʿܿ� � �$�6�H�Z�l�~ϐ� �ϴ���������X� � 2�D�V�h�zߌߞ߰� ������b�T���x��� ��d�v������� ������*�<�N�`� r�������������� &8J\n� ��� ���6�H� "4FXj|�� �����//0/ B/T/f/��x/�/�/�/ �/�/�/??,?>?P? �u?h?���?�? �?OO(O:OLO^OpO �O�O�O�O�O�O�O _ _$_�/H_Z_l_~_�_ �_�_�_�_�_�_o�? |?&o�?�?�?�o�o�o �o�o�o�o
.@ Rdv����� �>_��*�<�N�`� r���������oHo:o �^opo8�J�\�n��� ������ȟڟ���� "�4�F�X�j�|���� ��į֯�����0� B�T�f�x�ԏ����
� �.�����,�>�P� b�tφϘϪϼ����� ����(�:�Lߨ�p� �ߔߦ߸������� � �$�6ﲿ��N�ȿڿ 쿴���������� � 2�D�V�h�z������� ��������
f�.@ Rdv����� �>�p�b�+���` r������� //&/8/J/\/n/�/ �/�/�/�/�/�/? "?4?F?X?j?|?�?�? ��?�?2DVO0O BOTOfOxO�O�O�O�O �O�O�O__,_>_P_ b_t_�/�_�_�_�_�_ �_oo(o:oLo^o�? �?vo�?OO�o�o  $6HZl~� ������� � 2��_V�h�z������� ԏ���
�fo�o�o S��o�o��������П �����*�<�N�`� r���������̯ޯ:� ��&�8�J�\�n��� ������ȿ$���Z� l�~�F�X�j�|ώϠ� ������������0� B�T�f�xߊߜ����� ��������,�>�P� b�t��������*� <���(�:�L�^�p� ��������������  $6HZ��~� ������  2�����{���� ����
//./@/ R/d/v/�/�/�/�/�/ �/�/?b?<?N?`? r?�?�?�?�?�?�?�? LOO���nO�O �O�O�O�O�O�O�O_ "_4_F_X_j_|_�_�_ �_�_ ?�_�_oo0o BoTofoxo�o�o�o*O O�o@OROdO,>P bt������ ���(�:�L�^�p� ���_����ʏ܏� � �$�6�H�Z��o�o�o ���o؟���� � 2�D�V�h�z������� ¯ԯ���
��.��� @�d�v���������п �����t�=�0Ϫ� ��Ο�ϨϺ������� ��&�8�J�\�n߀� �ߤ߶�������H�� "�4�F�X�j�|��� ������R�D���h�z� ��T�f�x��������� ������,>P bt������ �(:L^p ������&�8� / /$/6/H/Z/l/~/�/ �/�/�/�/�/�/? ? 2?D?V?�h?�?�?�? �?�?�?�?
OO.O@O �eOXO����O�O �O�O__*_<_N_`_ r_�_�_�_�_�_�_�_ oop?8oJo\ono�o �o�o�o�o�o�o�ozO lO�O�O�O|�� �������0� B�T�f�x��������� ҏ.o����,�>�P� b�t�������8* �N`(�:�L�^�p� ��������ʯܯ� � �$�6�H�Z�l�~�ڏ ����ƿؿ���� � 2�D�V�h�ğ�π��� ������
��.�@� R�d�v߈ߚ߬߾��� ������*�<`� r����������� ��&��ϔ�>����� �Ϥ����������� "4FXj|�� �����V�0 BTfx���� �.�`�R�/v���P/ b/t/�/�/�/�/�/�/ �/??(?:?L?^?p? �?�?�?�?�?�? O O$O6OHOZOlO~O�O ��O�O"/4/F/_ _ 2_D_V_h_z_�_�_�_ �_�_�_�_
oo.o@o Rodo�?�o�o�o�o�o �o�o*<N�O �Of�O�O_��� ��&�8�J�\�n��� ������ȏڏ���� "�~oF�X�j�|����� ��ğ֟���V�z C���x��������� ү�����,�>�P� b�t���������ο*� ���(�:�L�^�p� �ϔϦϸ������J� \�n�6�H�Z�l�~ߐ� �ߴ���������� � 2�D�V�h�z��述� ��������
��.�@� R�d�v����ώ��� ,���*<N` r������� &8J��n� �������/ "/~�����k/�����/ �/�/�/�/�/??0? B?T?f?x?�?�?�?�? �?�?�?RO,O>OPO bOtO�O�O�O�O�O�O </_�Or/�/�/^_p_ �_�_�_�_�_�_�_ o o$o6oHoZolo~o�o �o�oO�o�o�o  2DVhz��_ _�0_B_T_�.�@� R�d�v���������Џ ����*�<�N�`� r��o������̟ޟ� ��&�8�J���� ��� �ȯگ���� "�4�F�X�j�|����� ��Ŀֿ�����z� 0�T�f�xϊϜϮ��� �������d�-� ߚ� �����ߘߪ߼����� ����(�:�L�^�p� ���������8� � �$�6�H�Z�l�~��� ������B�4���X�j� |�DVhz��� ����
.@ Rdv����� ��//*/</N/`/ r/�� ���/(�/ ??&?8?J?\?n?�? �?�?�?�?�?�?�?O "O4OFO�XO|O�O�O �O�O�O�O�O__0_ �/U_H_�/�/�/�_�_ �_�_�_oo,o>oPo boto�o�o�o�o�o�o �o`O(:L^p �������j_ \_��_�_�_l�~��� ����Ə؏���� � 2�D�V�h�z������� ���
��.�@� R�d�v������(�� �>�P��*�<�N�`� r���������̿޿� ��&�8�J�\�n�ʟ �Ϥ϶���������� "�4�F�Xߴ�}�p�� �����������0� B�T�f�x������ ��������,���P� b�t������������� ���߄�.�ߺ� �ߔ�����  $6HZl~� �����F�/ / 2/D/V/h/z/�/�/�/ �/PB?fx@? R?d?v?�?�?�?�?�? �?�?OO*O<ONO`O rO�O�O��O�O�O�O __&_8_J_\_n_�_��%�$SBR2 �1 5�P T�0 �  @?7 �_�_�_o o 2oDoVohozo�o�o�o �o�o�Q�o�_ 2 DVhz���� ����o��o@�R� d�v���������Џ� ���*��N�1�r� ��������̟ޟ�� �&�8�J�\�?���c� ����ȯگ����"� 4�F�X�j�|���q��� ��ֿ�����0�B� T�f�xϊϜϮ��ϣ�~�_�����!�3�E� W�i�{ߍߟ߱����� �������(�:�L�^� p�����������  �����H�Z�l�~� ��������������  2D(�:�z�� �����
. @RdvZ��� ���//*/</N/ `/r/�/�/�/��/�/ �/??&?8?J?\?n? �?�?�?�?�?�?�/�? O"O4OFOXOjO|O�O �O�O�O�O�O�O_�? 0_B_T_f_x_�_�_�_ �_�_�_�_oo,o>o "_boto�o�o�o�o�o �o�o(:L^ pTo������  ��$�6�H�Z�l�~� �����Ə؏����  �2�D�V�h�z����� ��������
��.� @�R�d�v��������� Я���؟�*�<�N� `�r���������̿޿ ���&�
�4�\�n� �ϒϤ϶��������� �"�4�F�X�<�|ߎ� �߲����������� 0�B�T�f�x��n߮� ����������,�>� P�b�t����������� ����(:L^ p������� ��$6HZl~ �������/  /D/V/h/z/�/�/ �/�/�/�/�/
??.? @?R?6/v?�?�?�?�? �?�?�?OO*O<ONO `OrOV?h?�O�O�O�O �O__&_8_J_\_n_ �_�_�_�O�O�_�_�_ o"o4oFoXojo|o�o �o�o�o�o�_�o 0BTfx��� ������o,�>� P�b�t���������Ώ �����(�:��^� p���������ʟܟ�  ��$�6�H�Z�l�P� ������Ưد����  �2�D�V�h�z����� ��¿Կ���
��.� @�R�d�vψϚϬϾ� �ϴ�����*�<�N� `�r߄ߖߨߺ����� �����&�8�J�\�n� ������������� �"���X�j�|��� ������������ 0BT8�J���� ����,> Pbt�j��� ��//(/:/L/^/ p/�/�/�/�/��/�/  ??$?6?H?Z?l?~? �?�?�?�?�?�?�/O  O2ODOVOhOzO�O�O �O�O�O�O�O
__ O @_R_d_v_�_�_�_�_ �_�_�_oo*o<oNo 2_ro�o�o�o�o�o�o �o&8J\n �do������ �"�4�F�X�j�|��� �����֏����� 0�B�T�f�x������� ��ҟ��ȏ��,�>� P�b�t���������ί ������:�L�^� p���������ʿܿ�  ��$�6��D�l�~� �Ϣϴ����������  �2�D�V�h�Lόߞ� ����������
��.� @�R�d�v���~߾� ��������*�<�N� `�r������������� ��&8J\n �������� ��"4FXj|� ������// 0/T/f/x/�/�/�/ �/�/�/�/??,?>? P?b?F/�?�?�?�?�? �?�?OO(O:OLO^O pO�Of?x?�O�O�O�O  __$_6_H_Z_l_~_ �_�_�_�O�O�_�_o  o2oDoVohozo�o�o �o�o�o�o�_�o. @Rdv���� ������o<�N� `�r���������̏ޏ ����&�8�J�.�n� ��������ȟڟ��� �"�4�F�X�j�|�`� ����į֯����� 0�B�T�f�x������� ��ҿ�����,�>� P�b�tφϘϪϼ��� ��Ŀ��(�:�L�^� p߂ߔߦ߸�������  ����6�H�Z�l�~� �������������  �2��(�h�z����� ����������
. @RdH�Z���� ���*<N `r��z��� �//&/8/J/\/n/ �/�/�/�/�/��/�/ ?"?4?F?X?j?|?�? �?�?�?�?�?�?�/O 0OBOTOfOxO�O�O�O �O�O�O�O__,_O P_b_t_�_�_�_�_�_ �_�_oo(o:oLo^o B_�o�o�o�o�o�o�o  $6HZl~ �to������  �2�D�V�h�z����� ������
��.� @�R�d�v��������� П�Ə؏�*�<�N� `�r���������̯ޯ �����
�J�\�n� ��������ȿڿ��� �"�4�F�*�T�|ώ� �ϲ����������� 0�B�T�f�x�\Ϝ߮� ����������,�>� P�b�t������� ������(�:�L�^� p���������������  $6HZl~ ������� ��2DVhz�� �����
//./ @/$d/v/�/�/�/�/ �/�/�/??*?<?N? `?r?V/�?�?�?�?�? �?OO&O8OJO\OnO �O�Ov?�?�O�O�O�O _"_4_F_X_j_|_�_ �_�_�_�O�O�_oo 0oBoTofoxo�o�o�o �o�o�o�o�_,> Pbt����� ����(�L�^� p���������ʏ܏�  ��$�6�H�Z�l�