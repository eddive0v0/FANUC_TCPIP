��   v	�A��*SYST�EM*��V8.3�0340 11�/9/2020 A   ����UI_CON�FIG_T  �� B$NUM�_MENUS � 9* NECT�CRECOVER�>CCOLOR_�CRR:EXTS�TAT��$TO�P>_IDXCMEM_LIMIR�$DBGLVL��POPUP_M�ASK�zA � $DUMMY�63�ODE�
4�CFOCA �5VCPS)C��g �HAN� � T�IMEOU�PI�PESIZE ޡ MWIN�PA�NEMAP�  �� � FAVB ?�� 
$HL�_�DIQ?� qEgLEMZ�UR� �l� Ss�$H�MI�RO+\~W ADONLY� }�TOUCH��PROOMMO�#?$�ALAR�< �FILVEW�	ENB=%%�fC 1"USER�:)FCTN:)WI��� I* _ED��l"V!_TITL�� 1"COOR{DF<#LOCK6%��$F%�!b"EBF�OR�? �"e&
�"�%�!BA�!j ?��"BG�%�!jI{NSR$IO}�7PM�X_PK}T�"IHELP� �MER�BLNK�C=ENAB�!? SIPMANUA�pL4"="�BEEY�?$�=&q!EDy#�M0IP0q!�JWD8�D7�DSB�� �GTB9I�:J�<BT_DEVICg1� &USTOM~0 t $} RT_SPID�r8DC@D*PAG� �?^C\ISCR�EuEF��UGN~�@$FLAG��@ #B�1  h� 	$PWD_A�CCES� E �8���C�!�%)$�LABE� $	Tz j�@�3
R�}	�CUSRVI >1  < `�Bp*�B� QPRI��m� t1^PTRI�P�"m�$$CL�A�@ ����Q��R��RtP\ S�I�}W � ���QIRT�s1}_�P'2 L3�hL3!x�R	 K,��?����QF�P�R�T�Q���S���P�!@<o��
 ���Q]o@oo�o�o�o�o�o Yo �o $6H�ol ~����U�� � �2�D�V��z��� ����ԏc���
�� .�@�R��v������� ��П�q���*�<� N�`��������̯ ޯm���&�8�J�\��n��PTPT�X������{� �s �{���$/�softpart�/genlink�?help=/m�d/tpmenu.dgp�
��.�@�r��&տ�pwd�� �ϟϱ���������� �/�A���e�w߉ߛ� �߿�N�`�����+�X=�O�����Q3`pb�b'b_� ($�߀���������������Q�Q�o|�z���$��k
y�p����e����  ��L"P����L�dz������P/`  1�b�����  �S)B� 1�XR �\�}!@wREG VED���0wholemod.htmD	�singlUd�oubltr�ip�brows�L�1��� �-?Qc��?Qdev.s�Zl��1�	t/����W/i/ {/E/�/�/�/�/�/?� �P(?:?L?^? p?�?�?�?�?�?�6�@ %?�?O�?0OBOTO#E 	??�O�O�O�O�O �O�O__)_;_M___ q_�_�_�_�_�_��_ �_oo/oAoSoeowo �o�o�o�o�o�o�o +=O?��� ������,�'O P�b�1�C�����aOsO Y�����:�5�G� Y���}�����ʟşן �����_?�9�g� y���������ӯ��� 	��-�?�Q�c�u��� ����y���
��.� @�R�d�vψσ��Ͼ� �ϟ���߽�Ϗ��N� I�[�mߖߑߣߵ��� ������&�!�3�E�n� i�{�I���������� ����/�A�S�e�w� �������������� տBTfx��� ������� Pb�+���� ����/:/5/G/ Y/�/}/�/�/�/�/�/ ���/�/?1?C?U?g? y?�?�?�?�?�?�?�? 	OO-O?OQOcO1�O �O�O�O�O�O
__._ @_;d_v_E_W_�_�_��Z�$UI_TO�PMENU 1��P�QR� 
d�QvA)�*default��OjM*lev�el0 *lK	 # o0cooao�sbtpio[23�]8tpst[1�huo�o�oCoUo =�
h58E01.�gif8	me�nu56y-pXq136zWr5zUt4]{Dq�������� *�uB�S�e�w��������<�prim=�Xqpage,1422,1������ #�5�@�Y�k�}��������B�Ȇclass,5�����'�49�D�М13@�v����������E�Ȍ53ڏ����0�B�E�Ȍ8�}������� ſD������1�C�nI�P�Qo{�*mm�`qkϥ�ϭfty�m<�o�amf[0�o��}	��c[164�g>�59�hq���{�Qx2�[}��qz}gw 5{�߹s[�m�F�X�j� |��ٿ���������� ���0�B�T�f�x����ϝ2�������� ��ڟOas�� &8d���� ϯ�14�^p����%�ȃainedis���//%/� �config�=single&>ȂwintpԀ0/ p/�/�/�/mJ�Qf´/ �/+e�/�o��?/?A? T?e?w?�?�?	?�?�? �?�?OO+O=OOO� qO�O�O�O�O�O�O%� _(_:_L_^_p_�O�_ �_�_�_�_�_}_ o$o 6oHoZolo~oo�o�o �o�o�o�o�o 2D Vhz	���� ��
��.�@�R�d� v��������Џ���]Nc�<��ϙ¿���iO���s�ͤ�ɟ�ϱ�u��|�f�؟>��4����Z����ߤ�6��u7���0�	�� -�?�Q���u������� ��Ͽ^����)�;�(M�_�>"41C�� �Ͻ��������)� ;�M�_��σߕߧ߹� ������2��%�7�I�[�m����6t���`������<$�74�� -�?�Q�c�u��,�����%	TPTX[2c09�,���24�0����Σ��18����P����0`2��`�1o�A�i�tv�������0�
�1��
ӯ�C:D$tre�eviewQ#�3��&dual=o�e81,26,4 ����~���/ /+/=/�a/s/�/�/ȩ/�/��;P�53 p��'?9?K?V/o? �?�?�?�?�?X?�?�?�O#O5OGO�/�/�1��/�2f��O�O�O �6hO�edit ���O�O,_>_P_��O �	_S\_�_�_�_�� �_oW�o�-o�So eowo�o�o�o�o�o?o �o+=Oat �㥝����� ��?B�T�f�x����� +���ҏ������� ,�P�b�t�������9� Ο�����(���L� ^�p�������5���ܯ � ��$�6�ůZ�l� ~�������C�ؿ��� � �2��_�_h�o�� �o�����������	� �-ߛ�9�c�u߈ߙ� �߽����ߣ�*�<� N�`�r��Ͽ����� �������&�8�J�\� n�������������� ����4FXj| ������ �0BTfx�� +����//� >/P/b/t/�/�/G�Y� �/}��/Y���?'?9? K?]?p?�?�??�?�? �?�? OO#O5OGO	� ~O�O�O�O�O�O�O5/ _ _2_D_V_h_�O�_ �_�_�_�_�_u_
oo .o@oRodovoo�o�o �o�o�o�o�o*< N`r���� ����&�8�J�\� n��������ȏڏ� ���/�/4��/X��?]O {�������ß՟��� g��/�A�S�e�x��� ����oO�����,� >���P�t��������� ο]����(�:�L� ۿpςϔϦϸ���Y� �� ��$�6�H�Z��� ~ߐߢߴ�����g��� � �2�D�V���h�� ���������u�
���.�@�R�d�� �*defaultq��B�*level�8˯%�ï������ �tpst[1�]��#y(tpio[23* �u(������	m�enu7.gif��
�13�	�5��
��
�4	u6 �
گOas��� �����//'/� K/]/o/�/�/�/�/F"�prim=�p�age,74,1��/�/??)?;?F"��&class,13@?v?�?�?�?�?M?_25�?�?OO0OBOE#T<�?|O�O�O�O�O�/�"18�/__ %_7_I_TO^26P_�_��_�_�_�_��$U�I_USERVI�EW 1"�"��R 
����_N�oo�m 8oaoso�o�o�oLo�o �o�o�o9K] o�,o���$� ��#�5��Y�k�}� ������V�׏���� ��,�>�P����� ����ӟv���	��-� ?��c�u�������V� `�ʯܯN� �)�;�M� _�q��������˿ݿ ����%�7�I���V� h�z�쿵��������� ��!�3�E�W�i�{�� �߱������ߒ���� ��S�e�w���>� �����������+�=� O�a�s��(������ ����'9��] o���H��� ���0B�} ����h��/ /1/C/�g/y/�/�/ �/Z�/�/�/R/?-? ??Q?c??�?�?�?�? �?r?�?OO)O;O�/ �?ZOlO�?�O�O�O�O �O_�O%_7_I_[_m_ _�_�_�_�_�_|X