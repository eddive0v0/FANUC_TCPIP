��   ��A��*SYST�EM*��V8.3�0340 11�/9/2020 A   ���	�BIN_CF�G_T   X� 	$ENTRI�ES  $QW0FP?NG1FU1O2F2OPz �?CNETG  ��DNSS* �8 7 ABLE�D? $IFAC�E_NUM? $�DBG_LEVE�L�OM_NAM�E !� FT�P_CTRL.{ @� LOG_8	��CMO>$D�NLD_FILT�ER�SUBDI�RCAP� H�O��NT. 4� H�9ADDR�TYP� A H� NGGTHOG��z �+LS/ D �$ROBOTI<G BPEER�� �MASK@MRUv~OMGDEVK�� RCM+ ;$�� �ިQSIZNTI�M$STAT�US_�?MAI�LSERV�  $�PLANT� <$�LIN�<$CLyU��f<$TOcoP$CC5&FR5&�JEC!�E�NB � ALA5R�B�TP�w#��V8 S��$VkAR)M�ONt&���t&APPLt&P�A� u%�s'POR� �_T!["ALE�RT5&2URL �}�#ATTA�C[0ERR_T7HRO�#US29��38� CH- �[4M�AX?WS_1;�y1MOD�z1�I� $y2 � (�y1PWD  ; L�Au00�NDq1T{RY�6DELA�3�z0��1ERSIS��!�2�RO�9CL�K�8M� ��0XM�L+ �#SGFRMn�#TCP�OU�#PING_RE�5�OP�!UF�#[A�C8�"u%_B_AUZ�@8��B�"COU!�_UMMY1�G2?��RDM*� /$DIS�� J@�Io/ 3 $A�RP�)_IPF�OW_��F_INFAD� ��HO_� INF�O��TELs# P~���� �WOR�1$ACCE� LV��RF:�!�ICE�0�Q�%  �$AS  �����Q��
���
�PV�1m@�W�  ���QI0AL�_�Q'�0 �X
���F��0���PBb;e���� #m��!�Qzo����$ETH_FLTgR  �Y.` �+ �������k��� #m2�kRSHA�R� 1#i # Pvo,8dX G|?�c��� ����B��f�)� ��M���q���䏧�� ˏ,��P��%���I� ��m�Ο��򟵟�(� �L��p�3���W��� {�ɯ��կ6��� Z��~�A�S���w�ؿ ������ ����V�� z�=Ϟ�a��υϻ���������@ߒgz _L��11�mx!1E.{�0I��z�1��>�255.�Ղ�&���@ey�2�ߒ�@�Ц߸�������3�߀��o��0�B�T���4 p������������5���_�� �2�D���6`�����������������6AM�Y�(MY���p��P� OQ� 8�<r ������%7 �Pgy�J �����	//-/���Cew/b,Q/���/�/�/�/�}�iRConnec�t: irc4//alerts�/ 9?K?]?o?5�/�?�?��?�?�?�?�0cP9a���?0OBOTO fOxO�O�O�O�O�O�O��O_�$�?3_�`( "_[_�/_�_�_�_�)���`a�i�R >j�U�Q�Qt)�eI �DMZcan�$T�CPIP[b�mXi(`=aEL`��ez�Q��`H!TB��o�rj3_�tpdb/ m�vQ!KCL�o�kv_|.��V!CRT�o��oF`�d!C�ONSG�j�as'monL�d