��   ��A��*SYST�EM*��V8.3�0340 11�/9/2020 A   ������DMR_S�HFERR_T �  $O�FFSET  � 	  /GR�P:� $�MA��R_DON�E  $OT�_MINUSJ � 	sPLzdC�OUNJ$REF,j�PO{���I$BCKLSH�_SIG�EA�CHMSTj�SsPC�
�MOVn �~ADAPT_I�NERJ FR�ICCOL_Pz,MGRAV��� HISID�SPk�HIFT�_7 O �N\m�MCH� S��ARM_PARA�O dcANG�o y2�CLD�E7�CALIB�Dn$GEA�R�2� RING,��<$]_d��REL3� 1�  	�FMS�V� +� M_LIF	��h(�t*���(DSTBl+_0z*_��=��f#�&WCL_TI}M
#PCCOM���FB� M� �M7AL_�ECI��P:!�%X{� $PS� �T�I��35�"L $�DTYk9�f1E�NDm4�`1�ACST1_4�22�93�9�4�95�96�6_O3VR�6� GA�7�2 �7�2�7�2�7�2�7�2��8FRMZ�6DE�DX�6CURLNHS�2sF�1�G �1�G�1�G�1�G�1�C�NA]1?(B0�$MΦ�PL� W ݀�STA:#TRGQ_M��k@KNVVSXZYZZY�I)ZI7ZIET �?VCMRPRU : � �B+_V:!�RHEP�T�SIZn�SDATvn �JOI� ��T��T��V��X�^�9P�(ORGlNEWl��T���T��V��U� �Yo  �$�1SS> O����a����}�`VERSI� ��g  ����aIRTUAqL�o�aS 1�h� ��� N �`��D/h O�w�����y �a��,��)�b�M� �q���������ˏG�����*�<�'�`����dP���������=gL�͸�ߟ?�����@� �%�7�I�[� m��������ǯٯ�>� �e�$��D��d  2x�u����� ����Ͽ������<d�A�S�e�wωϛ� �Ͽ�����������`5�(N�;�J�_�J߃� nߧߒߤ���������%��I�4�Y���$nS$ 1�lDj��E�� E�  �F@ F�5U��^���Z� 6!}�!}��,��� )�b�M���q������� ��� ��$HZ 揀eF����	�Ze�0� = C�,>P! ���i���/ �(/:/L///�/�/ �/e/�/�/�/ ?�/$? 6?H???~?�?�?a? �?�?�?�?�? O2ODO OOzO�O�O]O�O�O �O�O�O_._@_�O_ v_�_�_Y_�_�_�_�_ "Ҹ_o/oAo�_eowo �o�oZo�o�o�o�o�o +=�oas�� V������'��9�b,($1234567890]� o��[���������� �ُ����!�3�g� W�s�{�������͟՟ ���'�/�K�u�e� �������������� ��M�=�Y�a�s�������4 Ͽձ��P�LCL����� D??�  �+��N� ?r�]ϖρϺϥϷ���������8��VCoMRPR��2���dL�� ��0 +ߩ߻߂ߔ��ߔ�	� #�-��=�c�N��� ������