��  �A��*SYST�EM*��V8.3�0340 11�/9/2020 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  �  �ALRM_�RECOV� � � ALM"EN5B��&ON&! �MDG/ 0 �$DEBUG1PAI"dR$3AO� �TYPE �9!_�IF� ` �$ENABL@�$L� P d�#Uژ%Kx!MA�$iLI"�
� OG��f �%CAUSOd�!PPINFOE�Q/ �L A� �!�%/ H� �'�)EQU�IP 20N�AMr �72_O�VR�$VER�SI3 ��!COU�PLED� $�!PP_� CES( C p71s!Z3> ��! � $�SOFT�T_I�D{2TOTAL_�EQs $�0�0N�O�2U SPI_I�NDE]�5X{2S�CREEN_84no2SIGU0o?|�;�0PK_FI� �	$THKY�-GPANE�4 ~� DUMMY1d�TDd!_E4\A!R��!R�	 � �$TIT�!$I��N �Dd�Dd �DTs@�D5�F6�F7�F8�F9�G0�G�GZA��E�GrA�E�G1�G1
�G1�G1�G �@!�SBN_CF>"
� 8F CNV_J� ; �"�!_CMN�T�$FLAGyS]�CHEC��8 � ELLSET�UP � $�HOC0IO@� }%�SMACRO�ROREPR�X� D+`�0��R{�UHM�P�MN�B�! UT�OBACKU��0 �)DE7VIC�CTI:0�A� �0�#�/`B�S�$INTERVA�LO#ISP_UN9I�o`_DO^f7��iFR_F�0AI�NA���1+c�C�_WA�d'a�jOF�F__0N�DEL��hL� _aAqQbc?Yap.C?�Y`�A-E��#%sATB��d��AW{pT $DB� g"� =S�$MO�0B �0kq� \v� VE~a$FN!��pd�_�t�rdT_MP1_F�u2�w�1_~c�r~b!MO<� �cE D [�mp�a���REV��BIL0�!XI�� �R  �� OD�PT�$NOnPM��I�b�/"_�� m�蘁H��0DpS �p E RD_E�L�cq$FSSB�n&$CHKBD_YS�r�aAG G�"$SLOT_�H�2��� Vt�%��x�3 +a_EDIm   � �"���PS�`84%$�EP�1�1$OP��0�2qc�_OK8ʂ� e0P_C� c��+dR�U �PLACI4!�Q���( �a�p9M� <0$D������0pB�UOgB,�IG�ALLOW� �(K�"82�0VA�R��@�2B ����BL�0OU7� !,yq�`7��PS�`�0�M_O]d����CF�� X0G�R`0��M]qNF�LI����0UIR�E��$�wITCH^�sAX_N�PSs"�CF_LIM�t>=�SPEED�!����P��p�PJdV ���u�u3z`�P6��ELBOF� �W�@�W�p� ���3P�� FB���1��r�1��G� �>� WARNM�`dp܁�P���NST� �COR-PbFL{TR۵TRAT�P�T `� $ACC�Qa�N �r�pIأo"��RT�P_S\�r CHG@I�EZ�T���1�IE��T�Y1݀�� �x i#�Qʂ�H�DRBJ; #C��2���3��4��5��6*��7��8��9V3l�yM$�	3 @F TRQ��$�V����C�N�_U�pY�k�OpT <F ����𲨈#I2q�LLEC�7�"MULTI��b�"�A!cj DE�T_�R  4F STY�"b�=*�)2��o���pT |� �&$L�>��+��P��u�!TOt���E`�EXT����ၑB���"2(���Ӡt k0F�R�LƯ����� !D"�M��Qm� ���c0���"��G�1ćց�M���P��! q�Ջ��# L0�	���P �pA��$�JOB,�ǰR�0�TwRIG��$ d�� ������ �K� l���ļ�!C`�0b% et��F� CNG0A�qBA� ��x��
 �!v��� ��z�0�aP{`�R·&ΰ�f�Pt�a�!��"J�!�_R��rCJ�$�(J)�D�%C@Hӽ��z@h�P�4Z�@ '.�RO`�&̝סIT�c�NOM_�`���Sj��pT(�@�݉��1P�ǭ��RA�0��2&"�>�
$TF\V w�MD3�T���`UC1[�g�'�Hgb�s1q*E���\Ѐ�s�qŦgAŦsA�Y�NT�q�P|pDEeF�!)��G�PU8`/@�����AX���Ģ�eTAI~cBU�Fņ�|psQ* �� �'�PI�U)�P\7M[8Mh9�� k6F\7SIMQ�S)@KEE�3PATѠ"�%"�"$#�"~�L64FIXsQg+ ԭ�AdC_v�b���23�CCIh���5PCH�P�2ADD�6,AE,AG,A!H"�_�0�0_,@�f oA)�ԀzFK� '�=$#�"��4E��, l ���7zpF�CE�C!F+HS�EDIS�G�3��-�P��MARqG���r%�FAC
��rSLEW<����x;�M��MCY.����pJB����
a�C�Wv��U�V/ ��?�CHNS_E;MP��$GE gB݀_} ����pP�|!TC9f��y#a��� NdW#%I��r<��<��JR�И�SEGF�RoPIOj�ST�`�LIN׃�cPV����!�$0�����b�'��b�B��1` +`��	��a	` ���a�Pܠ��At��Py�QSIZ���ltKv�TVsE pz�y�aRS %Ѽ�uc@Q{k�|�`�x�Z`�`Ld�| `�vCRCɥ��!����t�`�%�9a˭9b��MIN@Q�9a7��q�D�YCk�Cz��le��50��p ��EV���F*ˁ_leF��N���P�Q۶�X%+4,���#0|!VSCAT�} AY��b1G"�2 �>�
/Ψ`_ rU@�+�w][��i %��7�k�R��3� �ߒ߱���5ġ�R�HANC��$cLG���*1$�0�ND�סAR�0N�K�a�q��acm�ME`�1��n�A0h�RA�Æm�AZ����X%O`�FCT���7`�rvS�P
ADI�O���u��pWP ��������Gv�BMP�d�p�D&ah��AESf@̓�W_NP�BAS���I9�4  �I�T�CSX@�w�m5��	$�1�)T��?sCb�Ny`�a~BP_HEIGH71���WID�0�aVTF�AC��u�!AQP80� �\�EXP+�L��@��CU�0MME�NU��6��TIT�1	�%��a�!�A1ERRL���7c \���q��OR�D���_IDG��QU�N_Od�0�$SCYS���4�ő�Iϡ�	�EVG#Ҍ�P�XWO����8���$SK�*2��T�(�TRL��9 ��� AC`�u䈠INMD� DJ�4 _Z�b*1K�*�W�PL�A��RWA.�tТSD��A�ת!�r@Y�U�MMY9�ª�10����¾��:	�A1P�R�q 
��PO9Sr��; ��[�$$�q�PLB��<�ߪS@��=��'�C�>4�'�EN5E�@T{�?S�S���RECOR.�@�H �O�@7;$L��<$��62�����`_q�b��_DL9�W0ROx@�aT[� ���b�.�F���������PAc���bETgURN�V�MR���U� ��CR��EWyM�bmAGNAL� �72$LA�e���=$P�>$P�٠= ?y�A<�C���@�DO�`������:���GO_AW� ��MO�a)�o����CSS_CNSwTCY�@A L� 0^�C`' ID[^�U2
2N��O����ـI�� B3 PNPRB^rzC�PIPOvI_#BY�R}�T�r���HNDG.�C �H�DQkSP�s*�SBLIO�F��0,��LS�D��0�N0�	FB��FE@��C��жE�cDO&a-sO�MC`@{�4�C�rH���WFPB�Q��SLA4�P�F�bIN� ��N3���G� $$���P]��v�@�v�ޕ���!o�"��#ID�&L�&9W�";$NTV*3"sVE 4��SKI���as�3�'2�b&aJ��&aM�mdSAFE�,d�'_SV��EX�CLU7ѻ���ONL`�#YcL����4��I_V8���PWPLYy�R��H[0�'3_M@�NPVORFY_S�2MSB�O@��k6�1�d~3�#Ot !5LS�EF��35�£1�`
%�P��$��t5�%�� Hy��TAx2�DP�� ��_SG� I � 
$CURB� _�
�B�������#H��3F��UNM��DZD@���l�{I`xA��J�F�EF��]IM�J @F]Bk��pOTb�k�ԋѠ�5�׿P�и@M� N�I��K��
RwPA�!(TDAY��LO�ADj��R�ӵ2 ��EF/�XILy��q}�OhPe�D��_RTRQ�QM !DF����P�r�S`<�ThU 2L�`���Qk�A���Q�Q'N 0�A�QA�t�RL���DUb���"җCAB�aO�B�N�S�QW`ID�`PWж��U/q� VjV_��P�P���DIAG��1�aP� 1$	Vb�HuTl��u�t� ��j���rRp�DQ�tVmE��Y@SW�a@d�p7`q��U�PM�pf�QOH�U�QPP�`&�sIR���rB��Fb �S��q��q�@3r��-x@ ��-uj#e�POwPx�P���uRQDWuMS���uA�u�b�tLIFEZ��C�p���rN�q�r�uxA�s��rI�xBCp����NC�Y��r�FL�AW�y@OV���vH�E'ArSUPPO$2���rS�_E�)E��_Xf�h���s�Zp�Wp�p�s���xA�ƙ�XZ����qY2�ˈC
�T�����eN�됕exAJ� v_ě�q��/���Q }`[ CACHE��3�SIZ�v*��"j�N� UFFIo�� �p���Ե3��6�����M����R �8�@KEYIMAG*�TM�ᄣ��D�謖�q���OCVsIE�`�S wP���Ll$@)#?� Q	��%���T�P�ST� !��`!���@!�VP!��0!�EMAILy�1Q��� __FAUL��U�8 �9��COUz ���T��|aV< �$��zS�PC`IT�#BUFF�)!F�O�y�o�D�B��nC�($����Ú�SAV �Ţ�`���`����|FP
�z���d� _0���"P_�OT������P[0�Ѓ� B��A�X��-�I���Wc7�_9G�s��YN_$q'�EW�RDuY��#rUMb�T��F+��fP^@D�&�X�0�����g�C_��&�AK��8�4B3��R��82�q��DSP���PCy�IM�pÖ��#�Æ`UM�:���K0d�IPm#�q	�o�CTH��=c�mPT���p�HSDIm�AB#SCz$��o�V� �`Я�&�`ӀQNV�!AGO�&ԑ�mƸ�F�a�аdR����,�SC8xbk(�MER4��FBCMP3�EiT�1�Y��FUX��DU���\���%2C�Df���z�u��R_�NOAUT�  Z�P4 �"U�IU�PS�C�@�C��1ϱב㍰��[/H *�L t� 3���֚@�0�#��� ���A��VQ��1�扑*��7��8��9���pT���1��1��1��U1��1��1��1��1 �2�2���2���2��2��2��2���2��2 �3�3��3���3��2����3��3��3 �4��_�XT�aQ\ <���I簉�p��3刡FDRxd/]T��V�0��p�r��rREM�`9F��rOVMI�>�AGTROVGD�T�gMXvINpG�fuaIND���r
��а$D�G��:sp��u�aD�VpRIV���roGEARI�IO�e	K7�tN�%(hQ�x�0h `��sZ_MCaMÀ�q;�UR��'^ ,�1?����� ?� �a?�!E�0�!�������_P}pP���`R�I�դ$�aUP2_� ` VPģTD����3�#?@�!�'�%ƻ��#BACܲaC T�Ţڠ�A);@OG.5%�CT����IFIq���x�:p�C5PTV�@�FM�R2
b 4�3LI��3 #/5/G/^|��u7%_���R_�A���`M�/-DGC{LFuDGDY_HLD�!�5�v��tRM���c���9? T�FS]��d P� �B�0��а$EX_�A�H�A�1kPl���@3[5�V�G:�
e �����SW�O�vD�EBUG4WR�eG�R� �U��BKUv��O1a� pPO�P�YoP��BUoP�MS�0OO���QS�M�0E�XPO���� _E f ��`���T�ERM�Ug�U �'ORIe0�Qh�Vz0GSM_80Ţ�Pi�U.��TAij�UU���UP�k� 9-��f$�Ua`�g$SEGfjx@E�LTOV�$US]E��NFI"��b�n �q+�d]dh$UFR02���a���f	@OT�gU�TA ���cNST`PA�T��?��bPTHJ� ���E�:��АbART+��e|�+�V��a�REL<z9�SHF�T�a q.x_SH"I�M^���f $`�r�xj)A�0OVR��NǲSHI_p&DU4�= %�AYLO��AֱI�ѻ# qk�%�k�ERV���q�yz� �g`<r4_0&���_0�RC�!9�ASYM	�9��aWJ�g��AE�#*qV���aUz�@`ֱ.u|���DuP��X�pYѪvOR`M�3&Z�GR�Q1Tl�oR��V�`�`A��B��m� �>�b671TO�C�a�QT!k�OP@Z2���}���303YOYߠREM�Rm�b9�Oѐ$�reT��R�e��h�Fq/4e$7PWR�IM���rsR_C�#tVIS`�sb�UD�#fsSV�W�B��b n� �$H.56�_ADDR�H�QGr2�'�� ��R��~�o H� S��Q�4_�`��_���_���SE�Al�HS��MN�A?p T���_����OL���v�x��ּPACRO��<�aS�ND_C���x�qٔZ�ROUP�Ӓ�_X���@��1 ��25���?�4 ?�<�@���?���?���2AMC�IO��W�D:��J���1Sq $� ;�_D� �PM����PRM_.�   �HTTP_��HQar (�OBcJE��"�/4$��LE�c��s � ���AB_��T�SS�S� �D�BGLV��KRL~ÙHITCOU�[BG��LOF�R�TEM�ī�xe�a7�f�SSQ ��JQUERY_FLA��G�HW��aQatZ����F�PUR�IO�h����u�у��ѿ� �IOLN�2u��
@C���$SL�2$INoPUT_�1$��bi�P m�D�SL��Qav��gߢԝ�=�s��=�H�E��F_AS:�Bw%0$L:0'ǈ:1�q��U`|p�a0Tժ�_��pHY� ������UOP�Ex `��>�����hᣐP�Ã�^���؏�x�1UJ	y �� � NE�wJsOG�g��DIS�3�J7���J8��7�!PI�a���7_L�AB�a3������A7PHI� Q��9�D�@J7J�� �@�_KEY {�K�LMONQa=z� $XR���~�WATCH_� ��s98��ELD.5y�� n�E{ ��aV8�(���CTR@s�����%R� LG�|����DSLG_SIZM�� &�@%,��%FD0I$; �Q2#�P=/" _� +��@��ЩR ��P��S��� �ťV>" ZIPDU�r��)N��3R}J���@P �A��]�d0U�-r�L6,DAUR�EA��/�h^GqH0��!��BOO2�~� C��ӐI�T�Ü>@��REC��SCRN����Dx��FR'�MARG�2 Ҡ�����N�"����	S3���W���A���JGMG'MNCHL����FNd�J&Kp'7PRGn)UF|(�pn|(FWD|(HL�)STP|*V|(e0|(,�|(RS�)H�+��C�t�#y���1P#'G9U籐$"'�r0&��d�"G`)WpPO�7��*��#M07FOC�wP(EX��TUIn%I�  #�2,#C 8#Cl p!�p��v3@����p�N�sANqA�҉b�pVAI��CLEAR�vDCS_HI\T�Bu�j�BO�HO�GSI�Gr�HS�H(IGN; ���Mm!��T٤�@DE�(4LL\�C���SBU�PR`���pmT4B$1EM��D����rRQa�����pW��Ρ4�OSU1zU2zU3zQYT�AR`� ����΁p�esԲs�IDX�	P�r��O�P��a�V+ST?�RiY��a� �$EfC kW��&f9f�V��V�� L���_�#�|p��U���וE��֕YU~�_ � ��� .�6���c �M�C � ���C�LDP?�J�TRQ�LI�[����i�dF�LG���`��srAD��w��LDutuORG��!21r��v�yxu��t���dд� ����t"5�du� P�T�`��bp�t�vRCLMC�t}��ẏ�YPMI����� Yd)�QRQ�����DSTBP��P [��h�AX�bi�k�>��EXCESy�7�R>�M��U���`O���dXQ>��V��Z�]�_AW�\�������:�`KB� \���n��$MB��LI��I�REQUIRE��cMON�
�a�DESBU��;�L�`MA�� ڰ ᛐ���Z�q;�ND>S�a�'��ړDC�2�:IN�7RSM�����@N���F3���PST� � �4}�LOC�VRI����UEX\�ANG��RY���� AQA��K�$t�1RBMF ��]���Y�b0�eǥ\C�SUP�eYP�FXS�IGG� � ����b�w� �c:6�d���%c��?��?�.���DASTACWk�E��E��t���N"R� t��+MD��I�)���@��-���Hp��ᥴX�<���ANSW!��(`Q�1��D��)����ܚ ��� ÀCU�; V� pY�YP��L�Oj�����5�W��3�E���U�MÇM�RR2B��� �(E�NA�q d�$CALIa��GtvA��29�RIN� ��<$R��SW0����)�ABC��D_J2SEu�Y����_J3��
��1S�P���Y�P���3P�"��Y�J�J�ChZ՞r�O!QIM��(�CSKPz��1$oC��Jq(�Q�ܺ�p�պհ�e�_AZ�r�V���ELQU��O�CMPs�)����R1T��G�1���5�F�P1�9�f�G�ZE�SMG0}��Օ`E)R�����PA �S�(���DI�)�JGκ`SCL����VE�L�aIN�b@��_�BL�@Y����Z�J�������䮀�IN�ACcR���	"(.��f`_u�!�<����<�܂�F���YP�DH��;����iP�$V����'A$@d�b��P`��qy��B��H �$B�EL��|�_ACCE�� �����OIRC_����pp�NT�Q�S$PS���bL��� (s��	1w@
PAT!H��_��_3..���_wQ�� ��rb��CC ��_MG !�$DD���`�FW�E�~���������D}E�PPABN6ROTSPEE��{Q�`��{QDEF�b���$USE)_��BCP��C�0BC�Y���q s�YN�A�A�}yм�}M�OU�NGRR� O8��Q�INC�m����h����i�ENCS��d�Y�&��f�# IN�RI.%���NT����NT2�3_U��`�A#LOWL�A~0��`�a&Da0Y�C���`�r��C,�(&MOS�@��MO�ǀ�wPE�RCH  ~#OV�� �'�Q�#F�d"&��F��
�gm �@w�A. 5LADw��v�)%p�d*_6z&TRK���QAYI�3쁏1.��5�3n������PMOM Bh��sp"�W������3azR��D�UЋS_BCKLSH_C.!E� �&� �-�?D�JJ���CLALBP'"�q8�0܀|ECHK�`�US�RTYJ�N����T:Seq}�_c�$_UM���IC�C�����C(LMT�_L wp� ṮWE]&P [P!U,�5A��+0gT8PC�!8H��`|���EC�p�bX�T���CN_��N����V�SF���)V g�a	'|�Q.
e�X7CAT�NSH���� ��eq
A
&F�/F��Z� PA�D�_P�E�3_�`���6� �a�3�d�EJG�p���c�O OG�W��TORQUY/Ւ#�9� ?�0�"��� r_W�5�4�C��<t��;u��;uI*C{IQ{I��F��.q�aҐxpѽ VC��0b�Z��r1�~���s��uJRK�|�r�v�KDB��M���M��_DL��:2GRV�Bt;���;����H_pL��b i�COSv��v�LN�p����� ��d���mq׊Ō�qb�Z���&�MY������TH��6�TH�ET0j%NK23���`��㣀CBe�C5B��C��AS���`mt����e�SB�󜶒p�GTS��(C��m�=�cM��ԃ$DU�@C7������ ���QF�s�$NE��ؠI���C)���T�AX�����h�s�s��LPHv�_�9%_�S �ңŅңԅ_����(����V��V���𪻬VʪV׫V�V��V�V�V�H���E�²��?aٸ׫H��H�H�H�H*�O��O��ONɹ�UOʪO׫O�O�UO�O�O�F_������Ņ�Ė�SPB?ALANCEQԃQ�LE͐H_X�SP��9�ņ9�ԆPFULC=�d�L�d�ԅ�&�1��UTO_<�@�eT1T2����2N�A��?�Ԗ��1�f�D�5���1TP0O�����,pINSEG��!REV�փ "!gDIFy5K�1�0�6��1�l0OB&�lA�E��72p?�A$�L�CHWARlA�B�a�5$MEC�H��%����FAX��1PJT��z���З� 
��q�%ROB� CR(2��R��MSK_����� P ��_WR ��r0�?{41	b4 �20�1#JD0���IN���MTCOM�_C�p��  �� 8�$NO�RE$#���t���7� 4�0GRr���FLA�$XY�Z_DA��nC DEBU�� ��t��� 0�$uCOD�[A ���2����0$BUFIN�DX2�C MO=R#�� H-��0 ���FB �0�JD$�����QVPTA�A+�2G6�� � $SIMUL�` 13�3�OBJE;ТAD�JUS�� AY_�I�A	8D�OUTp�`���0�_FI�=@T+p4  ��X�3p3�A�5�DrFRI(CXT&8ERO�` E3q[0��OPWO�p'��, SYSBU<q�( $SOP��A�U�3�PRUYNv��PAC�D���0_� NR�X��AB��PP� IMA�G[A-�G�P�IMY"$IN,��!#?RGOVRDM��� �P   #`W�L�_��an%�B�PRB�5PX�`QMC_E�D/ �� PPNq�Mx�"OQ@MY19NQ7 �M!SL;�'��� x $OV�SL��SDI{D�EX�S�&�SP1�"V3p�%N1q�03�78�"���M!_SsETp'� @�0�K2��AARI�� 
B^6_��j7�1v1�5� �P �<T����`ATUS@$TRCI�H%�3'BTM�7�1I��$�4NQ�3� '� DB-�E��"�2z�Ev��1!0l@�1EXE��0�A�!B*B�4S3��Z0.��0UP��9A9$Y�' XNN�7�qx�$�q�9 �PG���� $SU�B�1��1�1�3JM/PWAI,`P	3�E�LOP���$�RCVFAIL_CH��AR-�����Q�P�T�U�R_{PL�3DBTB�a��R�BWDV��UM�`TIG�( �ю4`TNL(`TjRR m���`
p	1XQ� �E�S�T�R�ADEF�SP�� � L�-���P_�P��SUCNI#�7�PmAR1@�&�3�_L�P�1%�Pw�&����`@�� "<0��)�T"NU�GKETb(p��`�P^R&� h� ARSIZE���1���naS� OR�3F�ORMAT��TTC�O� ja�EM����d�SUX�2G1P�LIOR&�  �$��P_SWIpu��!�1�cLLB&���� $BA̙`1�ON9AKPAM��0=y��BAJ5����2r68v��_KGNOW8cNrA�U9A"ߐDx� �PDC�ryPAY�[�t���y��wZ�sL�1��U!�PLCL_$� ! �s,qv�t�b"�vF�yCRP1O�z�2�tES���w�R4��w�tBASeE$�J�"W�_J�q
K�mA��fBu���r�qĮ�MA�X4P�`AL_ � $�Qh 1q�!���C[�D�sEfr�J�3����� T� P�DCK� ��T"CO_J3������
�hrl���� ���C_YQ>�  � �� �WD_1�z2�tD����n�^���m�|TI�A4��5��6[�MOMS ��ȓ��ȓ��B�@AD��억�\�PUB{R͔������f#��?` I$PI�$�Q M�=q�wk�B1�yk���0������iqRM�q�!Ħ~AĦ�A
��9�d5SPEED�G �b��E�T��T�EP -�C��Q+�Q�ESAM(�E����8�Ep{� m� $�� k�~@Ƕ�P_� ֹm�k�v{��ŵ��2,H��ǳIN̚� c��1���B�W�.�<W�w�GAMM��1>��$GET9" ��D;�u
��LI�BRcA�RI��$H�Ib@_=!�0k���E�h ��A����LW ��4�+��X��7���wP��CEUv�[ �0 7�I_b�x u��L�������ȓu���ٞ� �$^Ј 1���I�0R��D\��kAT��LEf�=q�1M�7��}��PMSWFLT]M��SCRsH7��`���!��~B�dSV&��P� A ������#S_SAqs$��eCNO;�C�1fB<� ����K�����S�C� ��hrǥ��m�D� a� ��� ���в�����U!C��������s ��dMJ�� � ���YLi�K���^SJ�|v!6O� K���BK�- ��O	W���9���M$P��p����DHc�"��1~B�`M��~T2� � $-΍$$W� �%ANG"�q� ���� !��5P&��o���(�c�#��X`O"����Zz�`�@� �y�OM��+�(�:�pL�^�p���CON@��eL;�_�B� | ၰ��ș@&��@& �࡚m'X&��.����e�$"���`X$$Pnma�PM0QU��� � 8#`QCsOU���QTHYPsHO/� HYS�`3ES-r� UE� ���S`O�d�   c$P�@�Ŋ2UN�0�b�@O��  � �P�p45�E��C�RROOGRA�1A2DO445IT�Ё1F0�INFO�� �%0g;�1AȬ!OI�2� (� SLEAQ���1��0k6F0yS�НD� 4#`�ENAB"20PTION�C�T̢/G�T�CGCFA� @b#`J$P��<2����RdH0OBG�2S�_ED�@  � ��{K�q�3��E�)�NU�G�HAUT<�ECOPY�qI0(�L���M��N�@�K^��PRUT �B�NV@OU�b$G�92DT�bRGADJ���bbX_ �R�$`pV�pVWnXP@nX[�pV�`Pz�N���_CYC"ZSN�SE�$ ��LGO����NYQ_FREQ0�Wb��a�d23L�p�b�PnQÓb���5CRE���#��I�F��s3NA��%�?d_G��STAT�U' ��*7MAIL䆲YsIN��$LAS�T�a���TELEM�A� �GFEASIA����H ��b�1���f;B����I �0���R=q�!� R�r�AB+A��Ex0�V@�a7vW�Cy��1�U8��I0�pd�lvRMS_TRs��@��s r7�z��akt� �T��/ 	�b 2� =�_+��ve� �w�r� �fe��c�NG�DOUa3;�NHC��RPR	 @��2G�RID�1+CBAR�S��TYCZROTIO㐾�³�&0_[d�!�P��B�OxD�� � �0�PO�Ra3��[���SRV�_`)˄ÆDI�T�^���������4���5��6��7��8�ぬ!F��A�#0$VALURs���d��"`�D�� E��u1��aa��=@#AN�㉒qaR�@a>��TOTAL��1���PW�SIJ���R�EGEN����#X�xxI3e%!��� TR^s0���_S��^����CVnQ�D��B8rE��cN��!��42�@ÓV_Hk�DA�~���GS_Y
�rfS��{AR�2� <RIG_SE�ch�Â2�e_80��C_v�`��ENHANC�!'� p�qEqb�Î��INT��� F<.3MASK��ipOVR�#P� N��@`a
�_�*6^�M��Bp[��f8��SLG��>��� \ ��e�H ���Sq�dDE�U��*7Ő�%�2�U�!�TEj  � (7��҆��J϶�"cIL_M`!d��P㈠�TQ� ��Ë1rpj�eV��CF��P_��op��M��[V1��V1��2�U2��3�3��4�4���ᄠ��������s��IN��VIB�� �İ����2��2���3��3��4��4 �ؾ���#"�������`%��׌ՠՌ�PLv`gTOR� ��INb�p�����  �p���MC_F� 	�B��L����B�ڐM�1IB���#� 1 ��)���KEEP__HNADD��!��$<p��C�_`�䂁��H ��O�!��P��p����G���REM���쑥�;�R�W�U�[de��HPWD w ��SBMo�*��G�1�2�� ~H COLLABu���a������ؑEb�0IT���0��7� ,� FLbq�$SYN��M�C��d�UP_�DLY��#2DE�LAJ �nbY� A�D�� QSK;IP�� Ļ�60aODD���t P_60 _2�g0^ ����	 	Q�	��	%��
2��
@?��
L��
Y��
9�QO�J2R�P��CEX]pT�SY��X�]P��Y�1�� RD�C��b�� ��@ReCg�R4ae��"d�ԇRGEr@sl�:�FcLG�!Pa�SW�IΨ�SPC�3�QUM�_Yt�2TH2N�&�# L 1�� �EF�@11�!� l�����C��AT4�ET1��7 s"k0o4j!�@Y�j!<3\�HOME�"�P<$2D"�J/\/n/�/�/�/�'3D"��/�/�/P�/?!?�'4D"�D?@V?h?z?�?�?�'5D"��?�?�?�?	OO�'6D"�>OPObOtO�O�O�'7D"ֻO�O�OP�O__�'8D"�8_@J_\_n_�_�_�%S��
�1�9 �q=#$��i�S�E��ٷ�a�LbݖJcIOq�rjiI�P��Į< �POWE��� �4` wGbה ���b$DSB��GNABqՔE C�) ���S232NPe� ���U�P�ICEUQrt�E|3 ��PARITá�ՑOPB��FLOW�TR`�c�3���CU+pM��U�XTn���U�ERF�ACtC�Uѐ�FbSCH�q� t�����_p��$L����OM۠9�A��T>���UPD�A$#�`T+`҃*�� 4�x�s!��FA�������RSPqpQ���� !�X$USaA ���Y�EXmp#IO6��pU�YE��b�_�ª�B�#q`�WRp��_�YD�����V?FRIEND���UFRAMδ��TwOOLȆMYH�����LENGTH_VTE��I���[��$SE�`��UFOINV_�@�5a�RGI���IT�I���XX�	�J�G2J�G1T�U�D�d�du���_Â#O_p@�py�ၻ��n�C	��zŔ�C ���ʖ ��G��zr2�� @ 9�qC���d�wu��ysF� ���p���X #�E_-M�pCT^�H��f�P�<u6�	�G#WV��z�G���Dh LOCK~�U� �������$� 2ߐ��~�D ��1���2*��2�3��3��� :����V��V=�"�=�
F�V��!Ѕ�/������p�xṿ�� ��Prƻ���������E������!��AC�PRs�!�b}�S���`��r<
��a� 0 5�"ؠ�V��ؠ���	�������
M�S��� ح�R�qda�¿$RUNN�`A)X2q��A��L�+"^��THICx� �w �u��FEREN�g���IF��x���I0����V��G1&�*�Є�1ٲ[�I�_J�FR�PR��
��R�V_DATA�q� RD�[ 
�A�L� �xՑ ��b{�  2� ��S��`�	ܧ �$ Z"G�ROU��!TOTܸ���DSP��JO�GLIYs�E_P�PrO��\7`��bv=K�p_MIR�.�2��MQ�O�APp���E<�o��t��SYS�E�ib��PG��BRqK���v$ AXIa  �⃃���Ҽ��A����H�BSOCd��T�N���16��$SV1�DE_�OPNsSFSPDO_OVR4 ����D� �OR+��PN��P,�F��,��OV��SFa���d�$�F�}�ja2㒓��ҁibL�CHH\RECOQV�n��WE�M�����RONs���_����� @�9�VsER��n�OFS9�C�Я�WDE���A����Rh��TRBq|6aY�E_FDOh�MB_CMkS B��BL��.�u��8āV摁��p��]�Gv��AM��i ������_M� [r�ec� T$CA��D:��HBK�q�vIO��,�a��PPA L1\D���bDVC_DB<���q�b���ja"�1���3���/ATIOi`jqcp��U�� �efCAB �����J���������__p�vSUBCPU�b�Sv��`_ ��p"�`'}���b"�?$HW_C� IpȺ��'ɣAx����$/UNIT��� � ATTRI���"��CYCL��NEC�A�Y�FLTR_2_FI#��h��fƂ�LP$���_S�CT��F_�'F_�,E2�*FS�a��"CHA��-7�1�Pr�2RSD  �b������a�`_T�PROX�MFpEM	`_��r��Ts2�� s2̍��5DI&��tRAOILAC���M��#LO�����5��ﰰ�����PR�S�̑{�dAC�p	���FUNC!��RIN됫�|�@�DEq3RA�@�� �C87`�CWARB�	#BLƑ�G�DA�K�!�H�HDA��AX�C�ELD�p�@S��2�A�@STI��`U��ѓ�$<�RIA��q�bAFQ P=���S��U ����3MsOI� PDF_�ؔ��qHpLM�FA�E�HRDY]�ORGEPH�0��|� P�UMULSE���`'*���0J(�JC�X��S�FAN_ALMsLVBs_aWRNfeHARD���v����p�@2$SHADOW��0��a�b��_`�+q�ї�_���vAU��Rx4\rTO_SBR��e���j� �|�A	sMPINF����!t6Q'sREGL���aDGBP��V�pL.�l�FL�%!���DAՀ_�P�C�M��N�Y�B�8V  ��� ]����$N�$Z�� ��Ҭ����� ��|�EG������qAR��#��2?��wP��AXE��ROB.��RED��WD���_F���SY��!���:h�Sr�WRIE��v� STR���`��7�E�!�����a���B����@CD� O�TO7q����AR�Y����.A���#�F�I��9�$LINQK�Q���y�_����6��8�XY�Z�bB�7P�OFF�
 �7�+��B��yB�����0}@��FI� ������yB
�_J��5������`Ȅҋ8��H�T�B�b�C0x�D�U �9AETURBa`XgSW���rX���FLz���#�p�u�Y���3\��� W1��K�M����31�DB`%��`'2ORQ�6�ѳC��}� DB��>��P��%����ќ\q:�OVEA���M 90=ѻs[��s[��rZ� �`X��aY�� X�O�~@ 91�P��B�F����=� S�B�_���s����SER�A	EBE��H� QC"�Aб������E�2��Q&QAX ���Q� �!�|�A ��+a�����@@��O����n������N���1 ����`��`��`�� `��`��`��`�� `��`�!��� �R�g�DEBU�#$��A�c�2��3�AB�GE�;�V�" 
�Ҷ���z!$� 
�$��$�@A$�O�$� n�$��$�N��T#��R\����LAB���� �GRO0��l� B_�1	ƞ�>� ���`�������a	�ANDàE ��<���aF� ��q��Z�0Qi�� ;�NTq`�cR�C�1=��
��~�p�SERVE��N�p� $q��@A�a!��PO�`X ������Q�p� � $��TRQ"m�
��Q�����R�2�oP@_ �� l=���fER)RҒ�IV����NgTOQ����L%�P�Ď�z�0G��%%��"��?�!P � �,��2 뺱RA~� 2� d�rD�  �p�$O��2�PvµO�CQ� �  >YCOUNT���FZN_CFG��G� 4� ^v2T�d �"���m W �F�s/� ��M�08b������X��0�FA~P���V�XA�������0���O A�P��b�pHELkpN�� 5ސB_wBAS�#RSR]v�m@;�S�!YQB 1T�B 2e*3e*4e*U5e*6e*7e*8�5!ROOGP� �:�3NL�q)�AB��@nC ACK�IN	T80�sU�``x1�)�_PUA��b�2OU��P�@^x"#�y0���b�TPFWD_KcARlfpZRE����PP�&Q�@QUE]zROB�2����`�aIb`�"#8�$C0Bv8�SEMա�6�`�A�STY4SO�0�dDI1�@r�1�aǿQ_TM�sMA�NRQAF8�END��d$KEYSWITCHS3h1#A�4�HE2�BEATM6�cPE�pLEks1����HUg3F�4h2S~(DDO_HOM�P�O�a� EF"�PR@���rS����v�@Oa<X �OV_M���`pPIOCM$��7����##HK�q� �D5�_w�U�b�2M��p�44�%�FORC�csWAR�R�9WO}M�p � @��T˓�`U��P�1�VU2�V3�V4��*Ox0L�R��^xOUNLO.0�dd�ED�a  �$�$CLASS `����.a-�-� �#`S�0+h�9`��?aIR�T?�,o>`AAVMގ�K 2 je� 0 � �55a�o�h\�o�m �l	�m-�k`��o2v7u�lV}b�ah����t{`BS4�� �1Li� <��� �2�D� V�h�z�������ԏ ���
��.�@�R�d� v���������П��� ��*�<�N�`�r��� ������̯ޯ��� &�8�J�\�n����������ȿڿ�����rCF`�AX�� `Ė�sl9�%�IN.��<Ŷ$�PR�0XEQ��}�`�_UPMIl��ja{`L�PR �ji`��tLMDG ��g�`��PIOF �k`d� �0�B�T�b�߅ߗ�x�߻���, 
� ��n��o�0�B�T�g��x�������yNG?TOL  �{�p�A   ��
�{`P�d�O �� @��=�O�a�s�6b�  ��u���2b�������� ����&J4Z���������� *<N`r�~�zPPLICA�1g ?je}�����Handl�ingTool �� 
V8.3�0P/58��?
88340��sF0!�755�����7DC3x�����ޝ��FRA� ;6*-  !�� GTIVqŵ>��#�UPn1 ��\�P>APGAPONf`�.�za� OUPLEDw 1�i� /0�3?E?W?�_CUR�EQ 1�k  P�a7a<�n�?�d�}��33b9b g���4H�5�22�:HTTHKY�?Kx�?�?ZO�?6O HOfOlO~O�O�O�O�O �O�O�OV_ _2_D_b_ h_z_�_�_�_�_�_�_ �_Roo.o@o^odovo �o�o�o�o�o�o�oN *<Z`r�� �����J��&� 8�V�\�n��������� ȏڏ�F��"�4�R� X�j�|�������ğ֟ �B���0�N�T�f� x���������ү�>� ��,�J�P�b�t��� ������ο�:��� (�F�L�^�pςϔϦ� ������6� ��$�B� H�Z�l�~ߐߢ��6s5�TO��/�#DO_CLEAN�/�$6��NM  �� a?�������g>DSPDRYR=�&p5HI� `�@q�8� J�\�n������������������m8MAX@�����17.X��-!*2-!�"PLUG�G0�*3�%PRC*��B^�b�'��O���
�SEGF� K���^�p�8J\n���LAP�(�3��� 
//./@/R/d/v/�/��/�/�#TOTAL�Py	�#USENU
"; �8?�2s0�RGDISPMM�C� o1C�@@I@
�"4O�5 �3_STRING� 1	�+
�kM� S�*
�1�_ITEM1�6  n�-�?�?�?�?�? OO'O9OKO]OoO�O��O�O�O�O�O�O�O�I/O SIG�NAL�5Tr�yout Mod�e�5Inp?PS�imulatedޒ1OutQ\�OVERR� =� 100�2In� cyclEU�1�Prog Abo�r[S�1;TSta�tus�3	Hea�rtbeat�7MH Faul�W�SAler�Y_ o o$o6oHoZolo~o�o�o �;�? �o�o);M_ q����������%�7��oWOR � �;o��oI������� ͏ߏ���'�9�K� ]�o���������ɟ۟�PO�;�Q��� ��6�H�Z�l�~����� ��Ưد���� �2��D�V�h�z����DEV���*���޿�� �&�8�J�\�nπϒ� �϶����������"�>4�PALT�m[� ��5߃ߕߧ߹����� ����%�7�I�[�m��������I�GRI3 �;��s���'�9� K�]�o����������� ������#5GYk��� R�m��} ���%7I [m��������/�PREG _�H �!/o/�/�/�/ �/�/�/�/�/?#?5? G?Y?k?}?�?�?�?]��$ARG_o�D ?	����1��  �	$V	[�
H]
G�W+I�0S�BN_CONFIOG 
�;IQHR�CACII_SA_VE  ThA�_B�0TCELLSETUP �:�%  OME_I�O]\%MOV�_H�@�O�OREP��_�:UTOBA�CK�ASM�FRA:\5+ �_5&�@'`�P�5'dX� q^ ,H5-�_�_�_�_8�_*o]T���0oXo jo|o�o�o�o5%Eo�o �o&8�o\n �����S�� �"�4�F��j�|���ࠏ��ď֏��  �PQ_3S_\ATB�CKCTL.TM�P XLED.GIF _$�6�H�Z���ZqsAkA0PIKNI^��U[E-S?MESSAGw@����A�0��ODE_D�@zFDV��O��ǟ-S�PAUS'� !�~�; ((O�2 �1��Q�?�u�c��� �������������;�I����TSK � 
�d__0PUP3DT����d��Ԗ�XWZD_ENB8��WJ��STA���1����1WSM_CFO@�5]E�7��GRP 2�} 	BB�  A����9XISI@UNT� 2j��C � �	z�� ���^ n�^ ��� %�� ��5*�����ϯ����π���0��T�W�i�M[ET� 2u�PN���J���^�SCRDV�1��P�EB��$�6�H�Z�l�~�]_5*Q{I����� ����(���L���p� ����������1�k��73QGRn����	��kNA�@�;	3Tn_ED��1˿
 �%-��EDT-���J��U /dD�@-3Sz5*�,B&o�Fs&  ��2�K� wʹ�E��	�-3�X5/|��/|/��k/�4 �/$/?H/��/H?�/�/7?�/5�?�/�? ?��?O[?m?O�?6LO�?�O�?�uO@�O'O9O�O]O7_ �Oe_�O�A_�_�O_�_)_8�_�1o��oxo�_�_go�_B9�o o�oDo���oD�o�o3�oCRS_���]���Ug��	 V NO�_DEL'GE?_UNUSE%�IGALLOW �19	��(�*SYSTEM*���	$SERVp*¯�Ȁ�REGх�$��ȀNUMx���	�PMUt�>��LAY�Я��PMPAL|��J�CYC10U��h�R�V���ULS�UH�
�j��ӃL���ݔBOXORI���CUR_ʐ	��PMCNVD��ʐ10~�0�T4D�LIȰß�ˋ$#MRߎ�&�&�ϲ ����̯ޯ���y	 �LAL_OUT �k��(WD_ABORo���m�ITR_RTN������m�NONST�OM �� ԸCE?_RIA_I�������˰F���U�c���_LI�M߂2` ԏ  N��Nϯ�<���m�`����  ?Ϡϲ��ϯ�
�����p��PARAMG�P 1U���Ύ�O�a�s�2�C>�  CV���f��z��ߵߗЇ�Б�Ж*�Р�Ъ�д�Ԛ�`����������C���_ǀ Cї��+�m��?�ɲHEC��ONFI�w�E�G�_P�1U� 49��������������E�KPAU�S�19� ,�uG�Y�C�}�g��� ������������1@U?e�!�M���NFO 1(�� �=����� ������A�/���%�q��w�Av���� Da���q~D�Q�6������ ˰O���ǩ��COLLECT_��(��pEN�`���\�INDE�x(���!��1234567890��������H,��)'/L/�| &/8/�/�{j/|/�/�/ �/�/?�/�/?e?0? B?T?�?x?�?�?�?�? �?�?=OOO,O�OPO@bOtO�O�O�"� �� ɶIO #"�����O_�a_s_�_WTR�2%#](�8Y
�O�^�P�$,]�Z��Y_�MOR"�%� � 9�Fe�Fi^oLo�opo �o�kb�#�&-mB򂦱?>�>����a�KTt�A�PM(���a�-=�Oa�s�ϗ�����^@�
����`w *c�PDBO�*���Ecpmi�dbg�C���U�:!����)�p/����S�  ��{be�-�̏��ܧ�a ��v����������g�^�)�=���fM���w���@ud1:˟���Z�?DEF )o7S�)ߑc�buf.txt��M� �p�_L64FIX +�Q���˓� د��ɯ��2�D�#� h�z�Y�������Կ��ſ
��.�f�x�_E ,� �l�~�`�Ϣϴ���p�IM�C�-�]��6��>̿��=L����M%C&c.�SdF�'�
%d/5ݤ`tձv���B!!� A*�B����B>BZA��,BA��A��;�B���DB�"C��<�C4�C�s��CC��D�2�FB�nE���E4��E���EC�2�y�bGɚ�g1�\D�y*T*�~**�}�Y�`U�x*�KCÇЯ��BDw�4  E	
��E�e�3Ec��E�t� F�3E?�ŚF�B� �F���F�Yf�F�% G�� �G	ڳH�3����  >�33� ;���a�v  �nf��q@�a5Y����b�pA�a�t�<#�eDQ�7���F��RSMOFST c'�f�G�T1#`uDZ�2!���Q,�*;�0�R�L��?���<�M^��TEST�0���FRz3SMx�C��A�z�*e�h��| C��B��3C�pn���*�:d�b2Iy4�<2T_�PR/OG ,k%^��/%PNUSER � �1��KE�Y_TBL  �-e1]�(��	
��� !"#$�%&'()*+,�-./�:;<=�>?@ABC�G�HIJKLMNO�PQRSTUVW�XYZ[\]^_�`abcdefg�hijklmno�pqrstuvw�xyz{|}~�������������������������������������������������������������������������������͓���������������������������������耇�����������������������A� LC�K#D#STA�Ti/0_AUTO�_DOG㺒�+IN�DT_ENB�/ a�"��/�&T2�/�6STOP�/�"S;XC� 25K�p�8
SONY �XC-56Q{�}�p�@���	�( АX5HR50�z-tx?�>y7�?�5Aff�:�O"O �?GOYO4O }O�OjO�O�O�O�O�O��O_1__U_g_�\T{RL� LETE6� �)T_SCR�EEN -jOkcs��PU0�MMENU 16� <O\�o �u�_oIo��&oLo�o \ono�o�o�o�o�o�o  9"oFX� |�����#�� �Y�0�B�h���x��� ׏���������U� ,�>���b�t������� П	����?��(�u� L�^����������ʯ ܯ)� ��8�q�H�Z� ��~���ݿ��ƿ�%� ���[�2�Dϑ�h�zπ���ϰ����b��S_?MANUAL"?�Q�DBCO� RIG��Ws)DBG_ER�RL� 7�[������ߴ��� O�NOUMLI I����dD
O�PXWO_RK 18����&�8�J�\�n�DBwTB_�Q 9<�����K,�D�B_AWAYW�^��GCP D=����_AL �/��SҡY!0�UD H�_q� +1:����0,R0�`T�PA�~���_M� �IS� ��@� ��OoNTIM�W�D�����
2#�M?OTNEND'"��RECORD 1�@� �����G�O�N<����z ���G��N r'9K���� ������#/ �G/�k/}/�/�// �/4/�/X/??1?C? �/g?�/�?�/�?�?�? �?T?	Ox?O�?QOcO uO�O�?�OO�O>O�O __)_�OM_8_F_�_�N�ex�_�_�_<_��_�_�_'o�N�U (o_oqo�_�o�o�o�o�NH�I�o�o�9$2o�N��� p��(�����N��_�K�]�����TOLEREN�C��B����L���O�CSS_CNSTCY 2A~�' h���Џޏ ����&�8�J�`�n� ��������ȟڟ�����"���DEVIC�E 2B~�  ��r���������ϯ�����)�����HN�DGD C~��Cz<���LS 2D\�;�����Ͽ�����=���PA?RAM E/����?�)���SLAV�E F~�J�_C�FG G/�)�d�MC:\��L�%04d.CSV�(��c����A &��CH��n�n�)�(�=�[��)�-�Z��j�X�W��JP����C�_CRC_O_UT H��<��+ϑ�SGN I�����\��18-MAR-25 08:16���)05��16�:01���� Ze�7-�)�)�*����o��Im���P�uG�=��V�ERSION ���V3.5�.20��EFLO�GIC 1J% 	��* �������PROG_E�NB����UL�S�� ,P��_A�CCLIM�����Ö7�WRSTJN����)���MO�
��x�INIT K%
��)� v�OPTp� �?	����
 	�R575)���7U4��6��7��5��
12���6��>��TO  ��@�t���V��DEXd��d��x��PAT�H ����A\���IAG_�GRP 2PI��|O�	 E7�� E?h D��� C� C ?��B���C��nk������C��Cm��B�N�BzoO�B�)�Bk��f383 �67890123�45���B� � A��A����A�A��O�A��A{�+As�Aj��RAbJAYc% x�@��ıp��G!��A�����B4h����x�
"����"��Q�A���A����A���A��� ��hAx~��Ao�7Af9X<��?$>��mF/X/е�h����("_��AY�;AS��TAM�^AGd�ZA@�A:�bA3%A+�-A$���)�/�/x��?�*@�;d�6����@{�@�u�-@o�@�i�7@cC�@\�j@V{N?\0�5?b?t?�??�@_��@Z^5�@T��@O��@IG�@C33�@<��@6�+;@/<@(�`J?\?��?�?O�8s� nE��@h�@b��!@\�0Vff@�Pt@Ihs@B��@;�bOtO�O �O�O�'6]^_p_N_�_ �_0_z_�_�_�_�_$o �_�_
olo~o\o�o�o >o�o��C"�!30�2xKA�@^>8Q�r��R?�  *u�^7�ŬFr'ş�5AFRu^@g�p�nv�@@�pp4pE�@[ Ah���u�C=+<���
=T��=�O�=��=�?<���<�p�q��xG� �?� ��C�  <(�]US� 4jr�D@�����"�A@w�?f�oX��mf��� �������ԏn��
���.�@��i?#�
b��\>�pn�^o��G���G�^@x���R����^8��ۑ�5甮�CnB�L]_u�T�&�P;�'f��d��aQ{���dD��  D�  C�����̯ޯ 8 ����V�ǯD�ïh�������3*Da��q�D��Q�7�f/´ �S�Կw������.���Rρ�!�'���t�>6��=���?�8xA��î�mYϧ� CT�_CONFIG �Q-��#��c�p�� STB_F_TTSd�
�����C�V����M�AU^����MSW�_CF��R-  �]z��OCVIEWf�SY�i���� �߽��������G�� .�@�R�d�v���� �����������*�<� N�`�r�����%����� ������8J\ n��!���� �"�FXj| ��/����/,/j�RCR�T�e&�!�,.V/�/z/�/�/��/�/�/�SBL_�FAULT U�I*n�1GPMSK���$7��TDIAG� V��e���1��UD1: 67�89012345�2��?�P�Ͻ?�?�? �?OO)O;OMO_OqO��O�O�O�O�O�O(� �>�;�
�?%_�ƟTRECPZ?l:
 z4l_?��?�_�_�_�_ �_�_oo0oBoTofo xo�o�o�o�o�o�O_�/_UMP_OP�TION��>*qT�RR���!9KuPM�E��>Y_TEM�P  È�33B�Пp�A�p�t�UNI7��şqF�Y�N_BRK W�Y�)8EMGDI_STA�u&��q ��p�NC�s1XY� ���o7�*�~y���d  ������Ǐُ��� �!�3�E�W�i�{��� ����ß՟����Xu "�4�F�X����f��� ����¯ԯ���
�� .�@�R�d�v������� ��п������%�7� I�[�u�ϑϣϵ��� �������!�3�E�W� i�{ߍߟ߱������� ����/�A�S�m�w� ������������ �+�=�O�a�s����� �������������' 9Ke�[���� ����#5G Yk}����� �/1/C/�o y/�/�/�/�/�/�/�/ 	??-???Q?c?u?�? �?�?�?�?�?�/O )O;OMOg/qO�O�O�O �O�O�O�O__%_7_ I_[_m__�_�_�_�_ �_�_Oo!o3oEo_O io{o�o�o�o�o�o�o �o/ASew �������_� �+�=�WoI�s����� ����͏ߏ���'� 9�K�]�o��������� ɟ۟���#�5�O� a�k�}�������ůׯ �����1�C�U�g� y���������ӿ��� 	��-�?�Y�c�uχ� �ϫϽ��������� )�;�M�_�q߃ߕߧ� ����E�����%�7� Q�[�m������� �������!�3�E�W� i�{������������� ��/I�Sew ������� +=Oas�� ������//'/ A7/]/o/�/�/�/�/ �/�/�/�/?#?5?G? Y?k?}?�?�?�?�?� ��?OO�?K/UOgO yO�O�O�O�O�O�O�O 	__-_?_Q_c_u_�_ �_�_�_�?�?�_oo )oCOMo_oqo�o�o�o �o�o�o�o%7 I[m���� �_���!�;oE�W� i�{�������ÏՏ� ����/�A�S�e�w� ������������� �3�%�O�a�s����� ����ͯ߯���'� 9�K�]�o��������� џÿ����+�=�G� Y�k�}Ϗϡϳ����� ������1�C�U�g� yߋߝ߯�ɿۿ���� 	��5�?�Q�c�u�� ������������ )�;�M�_�q������� !�������-�7 I[m���� ���!3EW i{������� �/%//A/S/e/w/ �/�/�/�/�/�/�/? ?+?=?O?a?s?�?�? �?��?�?�?O/O 9OKO]OoO�O�O�O�O �O�O�O�O_#_5_G_ Y_k_}_�_�_�?�?�_ �_�_�_'O1oCoUogo yo�o�o�o�o�o�o�o 	-?Qcu� ��_�_����o )�;�M�_�q������� ��ˏݏ���%�7� I�[�m�������ǟ ٟ����!�3�E�W� i�{�������ïկ� ����/�A�S�e�w� ��������ѿ���� �+�=�O�a�sυϗ� �ϻ���������'� 9�K�]�o߁ߓ߭��� ��������#�5�G� Y�k�}�������� ������1�C�U�g� y����߷��������� �-?Qcu� ������ );M_q����� ����	/%/7/ I/[/m//�/�/�/�/ �/�/�/?!?3?E?W? i?{?�?��?�?�?�? /OO/OAOSOeOwO �O�O�O�O�O�O�O_ _+_=_O_a_s_�_�? �_�_�_�_�?�_o'o 9oKo]ooo�o�o�o�o �o�o�o�o#5G�Yk}�_ �$E�NETMODE �1Y�U��  �P�P�U��{�pRROR�_PROG %³z%�V�&��uTA�BLE  �{�oe�w����w�rSE�V_NUM �r?  ��q����q_AUTO_ENB  �u�s�tw_NO΁ Z�{��q��  *�*�������Ā�+�*�<�N��HI�S���Q�p�_AL�M 1[�{ �2�T��P+O�˟@ݟ���%�S�_��.��  �{��r�j��pTCP_VE/R !�z!�5��$EXTLOG_7REQk��ቼ��SIZů��STK�������TOoL  �QDzs���A ��_BW�DJ��؆K�ԧ_D�I9� \�U���t�Q�rU�STE�Pa�s��p��OP_�DO��qFACTORY_TUNk��d̹DR_GRP� 1]�yށd 	�e�#��p�x������ �n�So� �k� ��� W��i�z�dϝψ��� ������	����?�*��c�N�@p�@���?���@%�:�j�
 F�5U҈�j��xd�����E7� E?p� D����L�D�>%��  C���K��B�  ;�  �A@E�o�@UUU�c�U��K��w>�]��>П���ѻ�{ E�F@ �����{�L���M���Jk�K��v�H�,�Hk{�{�?�  ��Q�9tQv+�8�?��6h�%7�{��]� p2J���1���/ �j g�,��FEATURE �^�UK��q�Handlin�gTool �� �roduCh�inese Di�ctionary���LOAD4�D St��ard���  NDIF�Analog �I/O��  d �- ��gle S�hift��F O�R��uto So�ftware U�pdate   �J70 mati�c BackupΦ�art Hgr�ound Ediyt���708\��_amera��F���D pr��nrR�ndImM��PC�VL��ommon� calib U}I q.pc��nf� Monit{or��wset��tr��Relia�b	 ��jp D�ata Acqu�is����� DiagnosD������ Docume�nt Viewe����
PC u�al Check Safety�� act.E�nhanced �UsGFrw ��\�weqpxt. oDIO � fi+� t\j7�en]dxErr� L*�  � �{s  $��r�� :����T "� FCTN_ Menu`v���t I�TP �In�fac% � 48\� G_ p� Mask Ex�ctg�� o��T� Proxy S�vH  5p��i�gh-SpexS�ki� " #1���#�mmuni�cC ons�apd�!ur ������"connecwt 2Pdin� �ncr stru�� I KAR�EL Cmd. �LE uaG"t\i�a�%Run-TiN�Env��"K��el +G sE S�/W�Li�cen��[GER�  �Book(System)��� R5� MACR�Os,x"/Offl� �Pa� MH��- �: \ac�1M�R� �)��Mec_hStopV!t�  ��0i���Mixx��E ��
� �0od
 wit;ch��Loa� �4z.�6 k G�1�3OptmUHM GGNW filG� HFz��g�' pmfO Multi-T= �i�4pa�PCM� fun�'{3M"PQo[�D QV�H�Regit0r�  � mpo� Priz@F�K _fcs �W g Num S�el�5��� DS� Adju� ���`W�
 4 S|Xtat�uQ/bUC�� �RDM Rob�ot��scove��� cctO Re�m�0�n���SS�ervH10@#CTX�PSNPX yb<2�� "K9$`�Libr���564@e�� �4H`ZU�SoY0t ssag�E�~� "�1�V�VLO�b/I- �pc
�`MIL;IB�mch1o Firm+�8� �b�"Acc` hXcT�PTX�;��� s Teln�0�m}B��5|��4Torqu
 imula�}�7Tou7@Pa51��Em�T_ �QC&V �ev. ocle�USB po,U � iP�a@Wd?USR EVxP+�Unexcep�tx�P�D{D{f}V�C�r�"�"�2�sV�D��j�cV�Hk u�ifoV�SP CgSUI�k��XC�6�X`Web Pl�V��9pjăa�+64.f��^ r>p�T�v�
J57À��vGrid�Qplay 76 (�X�`L&iR;�.��:K�\0ARC; 4 �120i��L#AsciiV!eRDAG�d��UplE@��� �@oCollW�Gu��� of^QޝPI  � 1�s� ��t�0tX8FK���Cy�p  2�*Porie  l�d�aFRL�1am�͉ RINT��M�I DevO0 (�&ax2 ,�0�%(}t�\rb�A/��Pa�sswo��:O"� 64MB DR;AM�

! 0ڢ�FRO�qG`��r�ciPvis�y6B�W�Welds c�ial�4 )��e�ll���!P�sh�K���wmrwd�c�XE|�( p�v� wmd�ty	 sPRa��PR0�t!1m@.)�8�D�P�����P+�D� 2b a���r�dr��Pb� q�DrT1�� eged� OL��Sup�r�AR8s�OPT "W� !� � d��; cro@�V  �SHe[�  ���
gq�<�uestZ;`LO SS��e�7tex E�$`�p$![b�UsCPP�@ �4YPVirt�W�St�e~�Pdp�n�x��  �� SWIMES7T f� F0���ui.�&���ĕߖ� аߕ�51s J����(Fr��Ε�II)�ߓ�on ��!���M!=��	QY�b��f>�t���mfV� �լ���Ҍr���? ���&P�3����8�b9���eie�߽�n\p���\R���ҭ`�A��2�p����!�
!����O����7 J5����5��8�1Q��\ar7���sXPR���k "��@}��b����`P���lnko����`1��RMJ����;���qM�����H54����j883]DER�N��Ffh�M/#el���չ1d/�� ����d0�/��|B�/��( �/��<��/��p�����.fd�/��AsSTC?��616�/��g HS|?z��as������1���?��0�?c�r W $O��!`��%rzP]O��t\awxOV4�` �O�$�a�O�ҵ��O�0���O��.EN _�D8�`<_��ite_?���v t_�� aO��IF{?�Ԉ`����) "s_�Epa��O-�>n1!Ot.IvTo5!�_��F���o^837�o*QogW-���o�/��X@�PDT4��_�ԓze�OHf4�_\7	9���MN������f�tro9?6�x�9i0���J59L��%����Ak��P����_p�o�Fp_-o0�@�?(�f1'?�pm_d��O���ٟ�O.�pe����m\�A��/_����'2.p�͆cW_��֮͠c�a/\ Ry8���(Las$����O_���0x���bo��<����I�̿"%� ���K��/?�siaf<Ϟd�?�NT+���Se����//`�C/�����'37��fiUf\����$SG���Ԁ6h��RDYaLS߱�oI�omw��_#�ps0����d�hVmj��93����E�ogW�P���ch\?�I��ퟓ� 8�o����rvi7�]�S�/������V(st�,��F���@�tl��u&5/����Td
�hWi��ݶSe��6O��sr��	��! ��y8P`��dr׏�o3PRI����a�O�/	X/��spr�ߕ��擇Li?/��3 H�6x/�d94'��6�3�q54 H�/v6353�/r4 H���&0�/�'��� X?v�72�Ie?�g13$;?��7�/58r?�'�6�/��Lo�_��t �ͅA�ϐOc�m�osK�!����O�����,�O9��O�OS�ua�lP_��8�?a_?�38�_��wr+��j83�?!�_]���NDSO-�f7O=�!��Y�ad�O9kl�o�s_#1�o��ip�#�-Et�op�RIN�,��/I���VA̳=SE_��0s
S���Z 0+ͅcmg�Z�� 4@�"�ut[/�of��`�M�r����@��N��596O_��4Џ"��U��#o(� I�c5%r_����e`���G�������c���AL"���lg303_U�oy� -<�t�
��	e�@t���RTU���h�z�xo���vo;��'O�52 ����4��'�Yu\�� vOA���4I`�FĿ
d -�ݕE���� (o�[�"qE3�yo��Wel_�p�������WMG���3aP@�Ϣ3wmg`[����߂�- ����On�45�?�fCM8k�IO��  �ߪ ������1���2�g�y�c R�;�Co���4(S�`�⯔�Ġ���3IF���� !�(�z�0at��N1T��q���R8��i5�᯳W2\��� O ��W?��˿ݿ￘��7��4SiZ/<���=�K�!�cl�i5\1sw/�S�AD���3CVt�Dt.�Q�mt�_�e���V�-aV�  /6��Nlo��D1��\�O�/C  �/�4 �/�i�e/��/1_�W62˟��o��/�eJ7��er9v�?�) "�?�svh�?
o�N� �?��.p[�tvhmoO�U749LOR`8r��OutlO?�t	\�?��j�_�//<�/h_ mpc��y�9\KO�j�_�/�_��uXP�/D�H8�gO}�oOnn�O�%N �߬u�'o���n]`�ߜ�oRCM�o�un@�_��$./_#���m  �H552�abe��q38BSR7�8�p�q�r0��libJ614�c�ATUP�@r�mc�p545zPs�gt�r6�V�CAM�3CR�I�p\rc�pCU�IF�  �q2�ptwd.f�NREN �rco�p631 � - Pr�pSC�HV� DiD�OCV>aIFL�C�SUJ18�0�p1�}�EIOC � ��4�p54�pR԰`4�9�pgm�SE�Tf�Sta�q�ql�ay,�p7�q�0�MASK�S�PRXYZaap��7f�C�pHOC�OC��3.3�r�p\�c΂51�p��qa�pp.�q39f�js50�q�ust3��LCH��A`
OPLG�1"�E��� "L3�MHCR�  08 (ĀSn@�Reg��CS�p��1H��p��q5�p0�8\�pMDSW o URGw�MD����sOP��\!�MPR�ra�4�Հ!�o��f��p! p��PC�M�H��R0БPath���p@aH�ՀRm����pTP���Հ�816�50�pgt��āS��ol,�99Ղ:�FRD�p(Qn�pMCN��cc�wH93�pLNP���SNBA@�rSH�LB��֑SMx�lrn?�63�p��q92�pL�HTC�pX�TMILVs�r�T���PAu�Y�sȡTmX>aEN��ELU��th��0�@`�8��qHѰr9��`ρ95Щp �Հ7��UE�V��adin(�C������pUFRI�e�eO�VCC�pt�VsCOY���VIP��'spd�[�I^�p��X͡tsπWEB��p��?�HTT�p �L2�R62�pCo�o?�CG��d�{IGt�
PRI���PGSN ng�I�RC��ne ��H�84�prd6�R7d��@�R��L�53�p�\lcl�q8�pDW" #4�6M� ��s52�8�R659�t�|�5�r dK�6��p��4�49�YpS���p5�̰L�06�pV�G MD�o�g, ƻ�66�p��ðAW�S�pJ643�LaIက�V��pzdҡ��u�GD����q�%�h�TY�� ���TQO�p<q�q6�g��p|� �-@��ORSY���R68�p3��O�Lp�ģOPIɰs{guK�SEND�$/аpLP�T�S��y���ETSɰ2!�6��U����-�43 m!D�VRu�ry:��IPN��onF�Gwene��oayt�D (S��E���I��0�֙���p�ytt\�sg��g "�ր�6h��L�yt\s�tr�ոA�ՀA��hk_t���yt����ces�լr��j7��mon.�՜A��d@�6��s-@�ׂ�yt4C6\�`Q���qh3��zDlli4�F�l1c�`�$rt{�� �¥���yt��w�x�U�vӐh8��nde��CAxV絰����N��zͰH��epen�戁�yt�T��Ģ��oqb3攢��h89��j��p��Pv�ed�����4 J7R80E5��0l��ձ`"t�644����� I�I���r�p����"�S��/л%��59�4G�tom���!�R J��� �֛Se3�ar3�E�t�32�%�Qsys�G�F ��������e;tr��urnk���f�20�x78���'�rn6������\jtET��
jo��ta.C����gr������� ����<���ge���01�7��2�yt�yt7�5b���Lj(���7. "P��T`dc��) ��	���0�r��1%at�@1O���p��daW(?��4tv/ 4oh��c8�}���s?yR�?�=losgm�?�;ild�?1<d�?N�@���0@$O�M���p1|O�;@x@���ytV��1���O_�	8�aic�C 2�9���C���7��6�E� �� `E?kedg?y=wm�`ORchl$_�2G&he>�4m_��7�5l�O 2�4O Oaw4OJmd9h\o�;dh2���oNsqz�o�kl���o�o��:��+F�e1t�'-�6J8"WQ��1 (F���pD1a�0��fr{F� x�� �f22.f�F;usS�pkg�M!�INgD�x���,���u��o�{��52�2�xsiRC�n� VM��^�992X�W� ��J9�b��st�'T��O 92\�6CMR/d#Z��O�;��ݎv'���tm�F����f8�vat��t+9>e��6sft"/��z_v(��ɟ?�4o��,�`��կK����vsw��8��Dni�o��lb ��蟮�����8W�\���vsmTڴaz�"����ο�"�of���ow�(�&��slw���f���`e�w�����*�vr�y4s�+N3GeN���Y�25:�oad��(�Na�NJ?��n�d�� "NwV  ;�(F8����rrd�6`��le &���C�U�4;��OFk7\��8���rk&�,��gl��P��g�Gt��il����~��   P�2^���38��r� ����0���J614��ATUPj���54�5����6F�V�CAM��CR�I!7� , UIFtB���2��ans���CNRE�'��63�1��RI��SCH��u65DOC�VN�ns� CSU��T|���0��HAoEIOC% "��54��R696{5\� ESET�W������7 C�u� MASK�t� 1PRXY�UJ N 7�ל�O�CO�om�513r�,,������ ��98\t����]�[�39�v!��oftwLCH!�g�OPLG:�950ai�P]P���e f,S�r��CS����g_lo��5� ��pDSW6�r7�0<!Pl DKO�PP4�PRQS#01� n Ad��\��X#PCMAa ¼�0�%���vd�v; �A
TX���0��1ADI�G� �!H ,S^�r723��9A�U�+ FRD!h#RwMCNr	H93���R2SNBA"�C�+ SHLB�	SM�p5�n m�J5�2�HTC���T7MIL6�Se����PO�0PA�86^*TPTX�VR�0{ELA4ool,�ԡ� P��8��\s�v���qSRVTf��95Q$95Aw\et� UEV��@a\AC!]�[AFR�!r��C!ol.�VCO��P��VIP�4e�� I6�t34[SX����WEB���@("�1T��,�l2tQ�, G�Eg\tkI�G�E#@`PPGS�"�PRC�4"TA�N��84��#R7��taQR�(
R�53�tRJ68���R66a5�2a- E��R6�5qr Im�5pa��l��573R64q���q5`MM� 061%�BFfx�R   ���WS!40�ACL�IQf9�PSniKaMS�E�Rn`���597{1TY�4776 J, TO��L����6�9 (k5�Pfer@ORS��CR68��\sun[!L%CSN� OPI1Tp�\0� ��Wsn.��L�E �bqS�fX�0ETS1T ����h#�0a�P �FVR� �,QN��4�GeneN�a
@�D�x���y�MG" �y���yg�_cc�y"�xcm�g_�y��yvth�yR�x3(�,�>�P��b��z1��z! cv�yon T�yh"�xhr�x�b݉1�`]�iA��y CV�yCP  �z��x��xt���	q��ypse������r;57� In���x�y͉576��(p�+�)� ����L� "yAl��w6\ab����j8<�B��h ���PR<�J8�zPcxC;�8�J�ps��9P��x96\{�(P��y�����A�xY`� �-��iv{�R DmM<�H7�zH6�{66�3�1�x�[�tor�������y�m�!��sZ�]�92����nalۺ�Й)�޸stK��}s3tr��ypsk���=�\p����xj932|�C��}�)��x8R�x2}�����.�|�޸_w���}hk�_k�FH��z9!�xk5e*�n�95
����yhe�z88�,�f�l.��H�eGt_w�y�"M�c� �� �zbak�H�Z�gent��h�\m���s���� ��d�� ���Y�;�(�Z�@�z
9Pf�yv�@��.��� ��� l�n�( l��gd��=
i��! xZ���+�00iB\��H[�H���� -�h�[�C" #��822��2�@}�OR��� ���iB/̿N@�"F���f��h@+�t=���tk� OR��ƈ�83�i1�t �˚�~nc+��fc䫚��5���835 �z����i�;�5:�B6�ri��ER���bv݉ (ˊng,�@�,4�*RȭY��k�xmo�`]/��p��+��ptp�z(�5�\pk�=O?�A�45 [ڈ��0�/�/ ?S�i�k߽�ij��
��?̚+�db��� s�50l�a��x���S��[d G�yϋ�c1e��0K�50�K�1�y�6h�Je��RDE��yqIn�t�
 Pa��(�9s\g{�H�919[ڸp�\:� Vi��tGool<?ވ	�J[��uppK/=_��vk {��K[��Z��Z��O �O�O�8�OK�H��?���_rj;*h�ndr�{�H]end��Ir�:�(�3��o>�73;���/�&7;*��{�X�j�|���"�4� � am_xO�v�e�ʘ���vI���oD�?|�xj{��� ��Tz{�] R5;�J9�;989ﭹ��(�_��p�m
�
�`�t���e�kR R�}�++R7�J L:;)C "���Kz�/p+z�x�d	�-�|�	�6{33�06 S�6I~R6�st�z���:�LND��IF �K�45��-con�{
C9�i�*ar �jyp�	�ds "X����ENl�y���s��l�gr��e-����856��`�z�rpi{�x=H�4� l�^�wj�! mr˛vv�:nn��}RC:| �� Jq9�Z����867��13J;6��8 �JT\�`��(iR��R|�"ٟc  �STD��.pLANG&�����r��ti����P��q���)0-�� E��k�g
��y` ��5<����R730��(�ޠ�8 (i��Er�rP��,�`��PCx��x���rvge��0����8���ge��a�<����	�.��is{io��ckin�� �R�(���pG�i� �����؁��j<	��PFK"��XAr��\@��BP4��!��d��aabbPbbb�����P�0�P��(1��SP��ޠ�FS J��J9]1��6859!	���02*4<627���Y���,����X���s\�GFSO�����sex��/�vr������&���RG�(R68'64�����#8	G (� CCR��I�v��cc�� "Ck�H���9�\RB�T}rgOPTN�4�4�2�4�?�?�O"Ocrg.8EF���8E��
DP�N��d�uDion= tEnd.tExaN�FINTtE��7tE�� ntEa�@tE�0"xtEHQtEhd\m�F�HD�F�uD\er!h�F���O�AitE��8sF�"UiretEh�uDtuDrh�GdCt�ed ������nG An�U�Y9p9�Ut2��8��0E���a�U�`t f�1���2��� m�U�a�U葠U-`As�U�ѠW
 ��1�ޭ��6h�U R�88�U851_f4<�`�Utiar�U����it� ��l"��M�R S�f`�fTX�P�U��epm�f"w #1�f! T�fy��fm�g��e�P�U� 2�U 70�Uon�jg���@_f J7r�Vipp�fon,�U����X�v4��j79b�fc��e]h98jg��"��\chp�WE�N�vd@Pb{StoD'�� E f�@�VgF0��el�gxѠU��jA8svY��f���6uh�arel�UKARNo�Comc�u�RĆeL*wp\ �V
+v�Y�u�fp\e�VA�N"���k�gpcp_f1a!I�[�f4y��wf
! Gf C�o�uarwf�FvІ84_f5 H�f�H84�v63 Hv�fH7�v779_fi24��7rw69*�+65�f1�g8p��V�75�VIC �f ;AP7v893���0R0���B�eck���Hs�
E����#fMNS+v�ПVՐ�V�P_f-]�_�Q�VX�\���tch믅ԠUw3\pSfWT"_f8dBe��Zhin_� ��03jgoX��(ROB�wOG���AUe@�A�^�HR�Pxf0lRuuyQuug_Sf̉�3uh523.�l=e*writy �6��2�6�5sv54�f�4І40����H�60�v0�h�[�08��+�=�O�a���18< ���68v�`��s�75^0��A�rw�7��h����וл�3z�v3Y� � �େ2f����� 29#f�p���\cib<f��;sbs�w��o scbP1oCjaa��Ly2%� -k��E"�74�9 wf c(W_�	`��XPF�&��wvF�E�X�Ϯ`�we�Vp��a\w�vTf͸�z50+�"#WV����֤u��2�tY �� ��nte�gx�����f04 (�g�x��D����BPX�k���I/��`o�d�@��G��pv k�F��ib�hp
om �wfE�A�f��Hfdn���z8Z�f��ؿ�ra�W�_�o�i �<�al�VVA�x�V�2�� 996�#fVCA��,�vast#/�q� ��"��dp/fyn:�fiL���58����D�Əodif��.e8D�P��q (d��o "���o��Rg�d9Ԑ�'G��strS���OsAW���wR73�v�16"� Rf�79r�2���iTra���c�h�/�wv"TqP+v̀��tpe�Mc�wor���+RC��59�8�� S5N+�809�?��C�fܸ"z\mߦ<�����RE��$F�L&0�pcz�6n�verv�gng_�N�746�_��S_�� Ch�?�� �]��8th��0�897i3�g�.��6�f!��y$��x���� T���;�&w& ����rk����`s�H�V�AGǧset�99�������$FEAT_AD�D ?	���Z�q�p��	x ������*�<� N�`�r���������̏ ޏ����&�8�J�\� n���������ȟڟ� ���"�4�F�X�j�|� ������į֯���� �0�B�T�f�x����� ����ҿ�����,� >�P�b�tφϘϪϼ� ��������(�:�L� ^�p߂ߔߦ߸����� �� ��$�6�H�Z�l� ~������������ � �2�D�V�h�z��� ������������
 .@Rdv��� ����*< N`r����� ��//&/8/J/\/ n/�/�/�/�/�/�/�/ �/?"?4?F?X?j?|?��?�?�tDEMO �^�y   x�=�?�?OO%O ROIO[O�OO�O�O�O �O�O�O__!_N_E_ W_�_{_�_�_�_�_�_ �_oooJoAoSo�o wo�o�o�o�o�o�o F=O|s� �������� B�9�K�x�o������� ҏɏۏ����>�5� G�t�k�}�����Οş ן����:�1�C�p� g�y�����ʯ��ӯ � ��	�6�-�?�l�c�u� ����ƿ��Ͽ���� 2�)�;�h�_�qϋϕ� �Ϲ��������.�%� 7�d�[�m߇ߑ߾ߵ� ��������*�!�3�`� W�i��������� ����&��/�\�S�e� ��������������� "+XOa{� ������ 'TK]w��� ����//#/P/ G/Y/s/}/�/�/�/�/ �/�/???L?C?U? o?y?�?�?�?�?�?�? O	OOHO?OQOkOuO �O�O�O�O�O�O__ _D_;_M_g_q_�_�_ �_�_�_�_
ooo@o 7oIocomo�o�o�o�o �o�o�o<3E _i������ ���8�/�A�[�e� ������ȏ��я���� �4�+�=�W�a����� ��ğ��͟����0� '�9�S�]��������� ��ɯ�����,�#�5� O�Y���}�������ſ ����(��1�K�U� ��yϋϸϯ������� ��$��-�G�Q�~�u� �ߴ߽߫������� � �)�C�M�z�q��� �����������%� ?�I�v�m�������� ������!;E ri{����� �7Ane w������/ //3/=/j/a/s/�/ �/�/�/�/�/??? /?9?f?]?o?�?�?�? �?�?�?O�?O+O5O bOYOkO�O�O�O�O�O �O_�O_'_1_^_U_ g_�_�_�_�_�_�_ o �_	o#o-oZoQoco�o �o�o�o�o�o�o�o )VM_��� �������%� R�I�[���������� Ǐ�����!�N�E� W���{�������ß� �����J�A�S��� w������������� ��F�=�O�|�s��� �������߿��� B�9�K�x�oρϮϥ� ����������>�5� G�t�k�}ߪߡ߳��� ������:�1�C�p� g�y���������� ��	�6�-�?�l�c�u� �������������� 2);h_q�� �����.% 7d[m���� ����*/!/3/`/ W/i/�/�/�/�/�/�/ �/�/&??/?\?S?e? �?�?�?�?�?�?�?�? "OO+OXOOOaO�O�O �O�O�O�O�O�O__ '_T_K_]_�_�_�_�_ �_�_�_�_oo#oPo GoYo�o}o�o�o�o�o �o�oLCU �y������ �	��H�?�Q�~�u� ��������׏��� �D�;�M�z�q����� ����ӟݟ
���@� 7�I�v�m�������� ϯٯ����<�3�E��r�i�{�����˽  ¸���� )�;�M�_�qσϕϧ� ����������%�7� I�[�m�ߑߣߵ��� �������!�3�E�W� i�{���������� ����/�A�S�e�w� �������������� +=Oas�� �����' 9K]o���� ����/#/5/G/ Y/k/}/�/�/�/�/�/ �/�/??1?C?U?g? y?�?�?�?�?�?�?�? 	OO-O?OQOcOuO�O �O�O�O�O�O�O__ )_;_M___q_�_�_�_ �_�_�_�_oo%o7o Io[omoo�o�o�o�o �o�o�o!3EW i{������ ���/�A�S�e�w� ��������я���� �+�=�O�a�s����� ����͟ߟ���'� 9�K�]�o��������� ɯۯ����#�5�G� Y�k�}�������ſ׿ �����1�C�U�g� yϋϝϯ��������� 	��-�?�Q�c�u߇� �߽߫��������� )�;�M�_�q���� ����������%�7� I�[�m���������� ������!3EW i{������ �/ASew �������/ /+/=/O/a/s/�/�/ �/�/�/�/�/??'? 9?K?]?o?�?�?�?�?>�9  �8�1 �?�?	OO-O?OQOcO uO�O�O�O�O�O�O�O __)_;_M___q_�_ �_�_�_�_�_�_oo %o7oIo[omoo�o�o �o�o�o�o�o!3 EWi{���� �����/�A�S� e�w���������я� ����+�=�O�a�s� ��������͟ߟ�� �'�9�K�]�o����� ����ɯۯ����#� 5�G�Y�k�}������� ſ׿�����1�C� U�g�yϋϝϯ����� ����	��-�?�Q�c� u߇ߙ߽߫������� ��)�;�M�_�q�� ������������ %�7�I�[�m������ ����������!3 EWi{���� ���/AS ew������ �//+/=/O/a/s/ �/�/�/�/�/�/�/? ?'?9?K?]?o?�?�? �?�?�?�?�?�?O#O 5OGOYOkO}O�O�O�O �O�O�O�O__1_C_ U_g_y_�_�_�_�_�_ �_�_	oo-o?oQoco uo�o�o�o�o�o�o�o );M_q� �������� %�7�I�[�m������ ��Ǐُ����!�3� E�W�i�{�������ß ՟�����/�A�S� e�w���������ѯ� ����+�=�O�a�s� ��������Ϳ߿�� �'�9�K�]�oρϓ� �Ϸ����������#� 5�G�Y�k�}ߏߡ߳� ����������1�C� U�g�y�������� ����	��-�?�Q�c� u��������������� );M_q� ������ %7I[m�� �����/!/3/ E/W/i/{/�/�/�/�/ �/�/�/??/?A?S?�e?w?�?�?�?�?�1�0�8�?�?OO1O COUOgOyO�O�O�O�O �O�O�O	__-_?_Q_ c_u_�_�_�_�_�_�_ �_oo)o;oMo_oqo �o�o�o�o�o�o�o %7I[m� �������!� 3�E�W�i�{������� ÏՏ�����/�A� S�e�w���������џ �����+�=�O�a� s���������ͯ߯� ��'�9�K�]�o��� ������ɿۿ���� #�5�G�Y�k�}Ϗϡ� ������������1� C�U�g�yߋߝ߯��� ������	��-�?�Q� c�u��������� ����)�;�M�_�q� �������������� %7I[m� ������! 3EWi{��� ����////A/ S/e/w/�/�/�/�/�/ �/�/??+?=?O?a? s?�?�?�?�?�?�?�? OO'O9OKO]OoO�O �O�O�O�O�O�O�O_ #_5_G_Y_k_}_�_�_ �_�_�_�_�_oo1o CoUogoyo�o�o�o�o �o�o�o	-?Q cu������ ���)�;�M�_�q� ��������ˏݏ�� �%�7�I�[�m���� ����ǟٟ����!� 3�E�W�i�{������� ïկ�����/�A� S�e�w���������ѹ��$FEAT_D�EMOIN  Vִ���ΰ�_INDEX������ILECOM�P _����7���-�S�ETUP2 `�7�A��  �N l�*�_AP2�BCK 1a7�  �)Ҹ�ϯ�%����ΰ:����� Ե��*߹�N���[߄� ߨ�7�����m��� &�8���\��߀��!� ��E���i������4� ��X�j��������� S���w���B�� f��s�+�O� ���>P�t ��9�]�� �(/�L/�p/�// �/5/�/�/k/ ?�/$? 6?�/Z?�/~??�?�? C?�?g?�?O�?2O�? VOhO�?�OO�O�OQO �OuO
_�O_@_�Od_ �O�_�_)_�_M_�_�_ �_o�_<oNo�_roo@�o%o�o�oF�z�P~�� 2��*.V1R�o�`* F`�cLpZepPCx|��`FR6:�"�~\��{T�� '��u�Q����w�Yf�*.F
���a	��s��Ռd�����STM �"�-��p��Y��`iPen�dant PanelY���HO���?����[�����GIF �6�A�"�ߟ񟆯��JPG����A���c�u�
��zJS�=��`�У+��%
Ja�vaScripti���CSZ���@����k� %Casc�ading St�yle Shee�ts�_`
ARGNAME.DT�
lD�\0��P�`��q��`�DISP*g�J�D����σ�����ϡ�	PANEL1��O�%D�8�x�k�}�+�2m���b���~ߐ�%�0�3��W�b� E����0�4u����b�����-�(�TP�EINS.XML�4���:\H���C�ustom To�olbar����PASSWORD��~}nFRS:\����� %Pass�word ConfigXoV��O ��o�?��u
 �.@�d�� )�M�q�/� </�`/r//�/%/�/ �/[/�//?�/�/J? �/n?�/g?�?3?�?W? �?�?�?"O�?FOXO�? |OO�O/OAO�OeO�O �O�O0_�OT_�Ox_�_ _�_=_�_�_s_o�_ ,o�_�_bo�_�ooo �oKo�ooo�o: �o^p�o�#�G Y�}���H�� l������1�ƏU�� ���� ���D�ӏ�z� 	���-���ԟc����� �.���R��v���� ��;�Я_�q����*� ��#�`�﯄������ I�޿m��ϣ�8�ǿ \������!϶�Eϯ� ��{�ߟ�4�F���j� �ώߠ�/���S���w� ����B���;�x�� ��+�����a����� ,���P���t����� 9���]�����(�� L^������ ��$FILE_D�GBCK 1a���� ��� ( �)
�SUMMARY.�DG�hMD:��0t Dia�g Summar�y1>

CONSLOG&	t��CConsol�e log�=	?TPACCN�/�%�4/?TP �Accounti�n�>
FR6:�IPKDMP.ZIPh/l
�/�/@�P Excepti�on�/n+MEMCHECK*/��@?�Memor?y DataA?��LN�)	FTAP��?'?�?K7��mment TB�D�?u7 >)�ETHERNET��?f�!OHOCE�thernet ~�figura�/�D�1DCSVRF�?�?�?�OQ1%��@ verify� all�O�M{,��EDIFF�Op�O�OO_R0%�HdiffQ_W�!�@CHGD1F_-_?_��_ f_�_S+�P�Y2�_�_�_Xo� �_ooGD3pNo5oGo�o no��fUPDAT�ES."piFORS:\ a}D�Updates �ListafPS�RBWLD.CM��hLr�c�P�S_ROBOWE�L�?<�aHAD�OW�o�o�of�Q3�Shadow C?hangesi���=�&�NOT�I�OA�S��O5N?otificqB���O�AJ?�n c��p���D��L�� 󟂟���;�M�ܟq�  �����6�˯Z��~� ��%���I�دm��� ��2�ǿٿh�����!� 3�¿W��{�
ψϱ� @���d���ߚ�/߾� S�e��ω�߭߿�N� ��r����=���a� �߅��&��J����� �����9�K���o��� ��"�����X���|� #��G��k}� 0��f��� ,U�y��> �b�	/�-/�Q/ c/��//�/:/�/�/ p/?�/)?;?�/_?�/ �?�?$?�?H?�?�?~? O�?7O�?DOmO�?�O  O�O�OVO�OzO_!_�OE_�Oi_{_�$FoILE_LpPR[p���_P�����XMDO?NLY 1a�UZP? 
 �
_�_ ._oR_o;o__o�_ �o�o$o�oHo�o�o~o �o7I�om�o�  ��V�z�!� �E��i�{�
���.� ÏՏd��������*� S��w������<�џ `������+���O�a� 🅯���8���߯�Z?VISBCK�X�Q>�S*.VD�0����FR:\��I�ON\DATA\��â��Vis�ion VD file\�j�����̯ ڿį�����4�ÿX� �|ώ�ϲ�A���e� w�ߛ�0�B���f��� ��ߛ���O���s�� ��>���b����� '����������� '�L���p������5����Y���}���$�ZM�R2_GRP 1�b�[�C4 w B� 	 �Q�k}h E�� E��  F@ Fǂ5U�/
h L����M��Jk��K�v�Hɿ,�Hk��?ǀ  �/h 9t�Qv8���6�h�%�A� � 3EBHeB��a `�E@i/�g��h @UUU�U��>�]��>П�;r8�	===E���<D�><��߳<�Ε�:��b�:/'79��W�9
@�8�?8�9��T/�Q/�/eE7� ?E?p D�D�/��D�  D� � Cζ/9
_CF�G c�[T ��/?0?B?�NO� �Z
F0�x1 }0�RM_C�HKTYP  B�P� �P�P�P��1{OM�0_MIN�0�
���0�PX��PSSB�#d�U�Pi�?	�3�O$O�UTP_DEOF_OW�P
�Y>?AIRCOM�0JO��$GENOVR/D_DO�6�RxL�THR�6 d�Ed�}D_ENBiO ^}@RAVCGe�7�� ��FnH� E�� Ga� H�� H�@Jh`�/O?_�G_X_{ ���AOU�@kN� {NB{8����_y_�_�_�_  C�� 	$o�XYoilCOmB��AVb~	��Y+O�@SMT�Cl��IZ �04d�$HO�STC�"1m��� 	
x&
{
:byeV�����z u� ��$�GH��p�	anonymousK�y��������� 	-�A�c� V�h�z������ԟ ����M�_�@�R�d� v���ˏݏ���� 7��*�<�N�`����� ������̿�!�3�� &�8�J�\ϟ���ïկ ׿��������"�4� w�X�j�|ߎߠ����� �������0�sυ� �ϩϫߜ��������� ���K�,�>�P�b��� s��ߪ��������� G�Y�k�L�p�� ����� $ 6YZ��~��� �	�-? /Su B/h/z/�/�/��/�/ �/�/
?-/_qR?d? v?�?�?��//? �?I/*O<ONO`OrO�/ �O�O�O�O�OO3?E?�&_8_J_\_n_�g�aE�NT 1n�i� � P!�O�_  �@�_�_�_o�_ +o�_Ooo[o6o�o�o lo�o�o�o�o�o9 �oo2�V�z �����5��Y� �}�@�v�����׏�� ������+��T�y� <���`�����埨�	� ̟ޟ?��c�&���J�QUICC0���p�!172.8?.9.225����A1���ү3���24�������!ROU�TER��`�r�ӿ!?PCJOGԿ���!192.168.0.10��~��CAMPRT$� �!�1�K�2ƃRT��O�a��ψTN�AME !�Z!�ROBO=���S_CFG 1m�Y� �A�uto-star�ted�4FTP�?[��?�O��O�� �������ߋO�(�:� L�o�]����������#��:4�F�X� 9�l��P��������� z�������#F��� Yk}����?�=�SM�65233)�
=_�,Rd v�K�����  %��5/G/Y/k/}/""q��?�? �?�/3?&?8?J? \?/�?�?�?�?�?�/ m?�?O"O4OFOXO�/ �/�/�/�?�O?�O�O __0_�?T_f_x_�_ �_�OA_�_�_�_oo ,ooO�O�OEo�_�o�O �o�o�o�o�o(: L^�o���� �� �CoUogoH�{ �o�������Ə�� ��� �2�U�׏U�z� ��������)�;� �O�q�R�d�v����� ]���Я����)����<�N�`�r�������_?ERR o�ʡ����PDUSIZ � 3�^L��ȴ�>�WRD ?�"���  ?guest-�!��3�E�W�i�{���SC�DMNGRP 2�p"�˰���3��-�K�� �	P01.05[ 8�� �����}> j  2��1�� � ����T���������������$���ϿQ�<�u�`�������  �  
���N(�P,�(����Q������[���l�� 8�#{�d�����"߾��_GROU��q*������	�����4S�QUPD  ��ȵX��TY������TTP�_AUTH 1r��� <!iP�endan�����8�g�!KAR�EL:*�����KC-�=�O�%�V�ISION SE!Tb�����!���� ��"� ��_6�H�l~��CTRL s�����3����FFF9E�3��FRS:DEFAULT�FANUC �Web Server����	�Ĵ�}�������W�R_CONFIGw t�� ���IDL_CPU�_PC*3�B���I  BH/%MI�N:,��M%GNR_�IO�����Ƿ1 N�PT_SIM_D�O&�+STAL�_SCRN& ���*TPMODNT�OL�'�+bRTY�(I!�&����ENB��'��-$OLNK 1u���Q?c?�u?�?�?�?�?52MA�STE~ ��52SL?AVE v��34>��O_CFG�?I�UO��OBCYC�LE>OD$_AS�G 1w����
 �?�O�O�O�O�O�O __1_C_U_g_y_�_\�;tBNUM�Ĺ=
BIPCH[O���@RTRY_CN *�"ĺB�!���P1��ȵ B;@Bx��>�Jo�1 SDT�_ISOLC  ���f��$J23_DS4�:��`?OBPROC?�%�JOG^�1y�;���d8�?��[�o�_?؟֟O|QNs��V����-�~o�h�`Y �A�_�bPOSRE��o�&KANJI_��0���/k�+�MONG zg��2�y� Ϗ����Ҿ)�0c	{,�9�T���e��_LY �R�_k�EY�LOGGIN@�����ȵ�$L�ANGUAGE Yk2$ 㑖��LG1b|�2����3�x�������O � '0,�� ��
q�3��MC:\RSCH�\00\��LN�_DISP }��?f�MKm�OCl�"@"Dzh#�A��OGBOOK ~K��w���w�w���X���-�?�Q�c��u���11����	 ���h�޿��������_BUFF 1@=���)� ����E�a�sϠϗ� �����������B� 9�K�]�oߜߓߥ�������DCS �>� =��͗�ֿ�M�l:�L�^�p���I�O 1�K No����������� ����%�9�I�[�m� ����������������@!3EY��Ex TMlnd���� ��0BTf x�������p//���SEV`�}��TYPln���/�/�/)-P�RS��P���bFL 1���`��?,?�>?P?b?t?�?�/TP袐loq"��NGN�AM�d��Ւ��UP�Su�GI�U\�e��1_LOAD�`G� %}�%DF�@GI6�?�[MA?XUALRM�Wk8�X\@�1_PR�T`�ԣ��Z@Cx���ꩦ��OV�9ŜC�`Pw 2��K �9��	q!P]  ��OQ�R9_$_6_ o_�]_�_�_�_�_�_ �_�_oo@oRo5ovo ao�o}o�o�o�o�o�o *N9rUg �������&� �J�-�?���k����� ȏڏ�����"��� X�C�|�g�������֟ ����ݟ�0��T�?� x���m�����ү��ǯ ��,��P�b�E����q���SGD_LDX�DISA�0�;��M�EMO_AP�0E� ?�;
  j ����*�<�N�`��rτ�Z@ISC 1��; �����T �A���ϛ�$��Hߙ��C_MSTR ��B-g�SCD 1����<߶�8����� ����"���X�C�|� g������������ �	�B�-�f�Q���u� ������������, <bM�q�� �����(L 7p[���� ��/�6/!/Z/E/ W/�/{/�/�/�/�/�/ �/?2??V?A?z?e?�?�?�?X�MKCF�G �vݽO�CL_TARM_�2��G�B P�2�@>OFD>{@METPU�C�@ۆ�~�ND�@AD�COL`E�@kNCM�NT�O tEo� �v��N5C.A�O�D�tEPOSCF�G��NPRPM�OYS�T@1��� 4=@��<#�
oQ�1 oU_�Wk_�_�_�_�_ �_�_o�_oOo1oCo �ogoyo�o�o�o�o�a�tASING_CH�K  �O$MODAQC��?���>~+uDEV 	���	MC:_|HS�IZEѽ���+uT�ASK %��%�$1234567�89 ��u)wTR_IG 1���l#E%��)����S�6�%CF�vYP�q>�At*s�EM_INF 1��#G �`)AT&FVg0E0`�׍)���E0V1&A3&�B1&D2&S0�&C1S0=ƍ)�ATZ׏+��H@/�W��K���A��@��j�ӟ����	� �� .�������;��� �Я⯕����*�<� #�`��%���I�[�m� ޿鯣��K�8���� n�)ϒ�y϶���{��� ����ÿտF���jߡ� {ߠ�S���������� �����T���+ߜ� ��a���	�����,� ��P�7�t���9��]� o�����(:q� ^��=�����XNITOR�@G� ?s{   	?EXEC1�3U2%3%4%5%T�p'7%8%9�3 ��$�0� <�H�T�`�@l�x���2�U2�2�2�2�U2�2�2�2�U2�3�3�30�+qR_GRP_S�V 1��� (��a��\��*X�>�<���A����#c>��~Z}�q_D{�~�1�PL_NAME �!#E0�!�Default �Personal�ity (fro�m FD) �4R�R2�! 1�L?68L@�1P
d d�?v?�?�? �?�?�?�?�?OO*O <ONO`OrO�O�O�O�O�O�OJx2e?_ _2_ D_V_h_z_�_�_�_r<�O�_�_�_o"o4o FoXojo|o�o�o�i�V��_�n
�o�oNtP �o*<N`r�� �������&� 8�n��������� ȏڏ����"�4�F� X�j�|�K�]���ğ֟ �����0�B�T�f��x���������Ү �FnH F��� G=��'�   #�����"d��� 0�B�&�d�r��׭Ҫ�\�������ݿ� ͸��� ��0�6πT�vϿ �ϩ�ͰA�  ��˿��Ǹ ]0���ƿ3�¿W�B�@{ߍ�x߱�B5K3�9�^0`�!0 �� �0�� @oD�  ��?�����?� ��!A������$��(;�	�l�	 ��p�V� ]0�M� � � � ��l�r� K(���K(�K ���J�n�J�^_J&Ǔ�2�������� @Y�,�@Cz@I��@�������N�����f����_�I���S�Ѭ�Ä��  �<��% �3�������!?s8y��
�/�!�x����T� ܌��������}��  �  �������  ����������	'� �� 0I� ?�  ������:�ÈTÈ=����l��	�(�|�����Ѧ����ψ��N@0�  �'���@2�?�@���@!��૑@)��C@0C���\CI�CM�C:Q�� ��ģ�%%��_�� ��B��0�@0��l@� ��!Dz���V�//�+/Q/���� ��H@q)q�%  ���+��� p�!?�ff���/�/�V/ ���/;��8 � !?/:��D4�� \6Pf8�)c�\�\���?Lv �$��;�C�d;�pf<���<��.<p���<�?L:��ݧA����d����?offf?�?&@ސ�@�� B�N�@T�,E�	�� 	A���dO�O�7 H��/�O�O�O�O _�O $__H_Z_E_~_�MEF�m_�_i_�_UO��_yI�_2o�XC��E���"Gd G;ML!o�omo�o�o�o �o�o�o�o$H�� iww9��_�o�@U��*�<�ڪ��� �/�6������ď��菎�A�A���ł�C؏=�ԏ��X���񨑟,�����  G�P��"@�<��E� C���s���x�؄�(�����/�B��/B"�}A���#A��9@�dZ?vȴ,���~��<)��+� =�G���j���q����
AC
=C������년� ���p�Cc��¥�B=����ff�{�,�I���HD-��H�d@I�^�F8$ D;ޓ�ܪ�̠Jj���I�G��FP<���QpJ�nPH�?�I��q�F.� D��Ɵg�R���v��� �����п	���-�� Q�<�Nχ�rϫϖ��� �������)��M�8� q�\ߕ߀߹ߤ߶��� �����7�"�[�F�k� ��|����������� !���W�B�{�f��� ������������ A,eP�t�� ����+; aL�p�����=(����3:��1���%�3�V�8�/"�(/:/�!4M��T/f/F1ϴ=Ӏ/�/4U?e'��T9�-�)��/�/?�/4?"<]�P�2Pf>�q��?���?�?�?�?�9���(�?�?/OO?OeOPO�QB�hOzO�O�O�O �O�O�?t.__R_@[/X_b_�_�_�_�_�_�Q{f�_�_o
o�@o.odorj  2 �FnH"�F��"�G=��B# ��#C9)��@|�@��o� �q�o{E�� �F��`�H C�����oA`��kE�0wGa�O�����{?ސ�q �\dR  zq `�
 �!�3�E�W� i�{�������ÏՏ�p������q ��P+��~Y��$MS�KCFMAP  ��%� �^f�q�qp�D�ON�REL  X5�[��0D�EXCFENB��
Y�����FNC����JOG_OVLIM��d�����dD�KEY��z���_PAN�����D�RUN����>�SFSPDT�Yw0������SIG�N����T1MOT�럜�D�_CE_�GRP 1��%[�\�O��O�&� �d�Q��u�,�j��� b�Ͽ��Ŀϼ�)�;� �_�σϕ�LϹ�p� ���Ϧ��%��I� ��m��fߣ�OvD�QZ_EDIT��U���TCOM_CFG 1�Q������"�
��_ARC_�X5ؙT_MN�_MODE������UAP_CPL�F４NOCHEC�K ?Q� W5�H��������� �'�9�K�]�o�����������v�NO_WAIT_L���׾��NT���Q��{�_ERRȡ2�Q��1� ��t���H*�����`��OI�Px 	��K��!8��?0|4�pBP�ARAMJ�Q���	��7so�� =�`345678901�/ *� ?/Q/-/]/�/�/u/�/�/�+�7�?<��7?��UM_RSPACEN�'2$�p?z4��$ODRDSP�E㌦��OFFSET_CAR�Ќ�6�DIS�?�2PEN_FILE�0�$���֌1PTION_�IO
�=�@M_P�RG %\:%$�*IO[N�3WORK� �Χ�� ����F7��Bh��� ��d�@(7�A	� ��x�A5��c���0RG_DSBL'  \5���|_��1RIENTTO��9�C��pZ��a��0UT_SIM_EDGX�+��0V�0?LCT �%��x�Dx=gT_PEXh���?�TRATh� d��T�0UP )�u^�Ӡ�ooX�_:oHi�$�2ǣ��L68L@}�_S
d d'? �o�o�o�o�o�o�o 1CUgy��@�����I2~o '�9�K�]�o���������ɏ9�<���� )�;�M�_�q������� ��H�j3�H1`��XRP�C�U�g�y� ��������ӯ���	� �-�?�Q� �2����� ����Ͽ����)� ;�M�_�qσϕ�d�v� ��������%�7�I� [�m�ߑߣߵ�����X�ϡ��*��S�H�Z�?�}����@��&?������� �����+�I�O�m�����?@����� A�  ������� ���M8q\�����z�d`O�P1��k����sd`�R0 ���D$@ @D�C  DD?Q�D	��U� � ;�	l1	 ���p�s& ' j � _� � ʉ��� H<zH<W��H3k7G��CG���G9|�+c	�H
��� CC9P/9P49S;Q9�/��9  ���  1!�H7 3�����/1/C/�BY����XQ��^�H�<Pq/ ܩ/�"2�#�3�.��    ��0�� �  0�6�/?�	'� � M2�I� �  ����
=���0q?�;�#&�(�3�/ ��A�?4;�B�?r�NEPO  'VP�3D�b CEPC��+\Cf Cj Cn/@O|ROߑ  ���~�D%%���� �B`���FEP�E˜@XP�E5z�_s/8_#_�H_n_�"�� ��H]2�Y�A�U  ��C�H�A�0p�Q?�ff���_�_�s_ ��o(k�18 �0>oLj-�!adTW�0yfP�h�Y�yy�3�?L�0�T�!;�C�d;�pf<���<��.<p���<�?ij��WA��Eل1d�31��?offf?�@?&+p�VT@��=r�N�@T�IuՉ�� &q-�0!��w e o������ A�,�e�w�b������� я����l���O���CE���2Gd G;�|>��� ��ß���ҟ���� A�,�e�����V��� �د6���r�#�5�G�Y��Z� �_�f���@����̿��A @!A�@%���5�C��Z�x��/i�?�؈�p���ϳ�U�P��2�]!YNE� CU%�̣�Ŀ����E��@I�!t�B�/�B"�}A���#A��9@�d�Z?vȖ+~��~���<)�+?� =�G�(߇����q���
A�C
=C������녡� ���p�Cc�¥��B=��ؿff�{��I����HD-�H��d@I�^�F�8$ D;���ڭ�̠Jj��I��G�FP�<��QpJn�PH�?�I�q�F.� D��E �τ�o�������� ���&��J�5�n�Y� k������������� �� F1jU�y ������0 T?xc��� ����//>/)/ ;/t/_/�/�/�/�/�/ �/�/??:?%?^?I? �?m?�?�?�?�?�? O �?$OOHO3OXO~OiO@�O�O�O�O�O��(}�ϳ�3:�O�a��<)U�E3�V�_+_�9R�E_W_t�4�M��q_�_t��=�ӝ_�_4Ue'��T9�]�Y	o�_�-ooQo?lz�P�bP�n�����o�O�o�ox�o�i���(�L7\�mt�B����������o��K�9�o�]�/ u������ŏ�ُ�{f��9�'�]�K������  2 F�nH��F�Щ�G�=��B@P!�.�C9F��p��@2���	��~C�E�� F����H C���S�b����������¯Dԯ��?����y��C�C�|�C�}�
 ۯ>�P�b� t���������ο�����(ϧ�� ���m[�~Y��$P�ARAM_MEN�U ?�U��  �DEFPULSE�4�	WAITT�MOUT��RC�V�� SHE�LL_WRK.$�CUR_STYLv����OPT�N��PTB����C��R_DECSN�� teG�A�S�eߎ߉ߛ� ������������+��=�f�a�SSREL?_ID  �U�a��u�USE_PR_OG %p�%b���v�CCR����a�x���_HOST !p�!�����AT�`��8����:�|t���_TIME������a�GDEB�UG��p�v�GINP_FLMSK�����TR����PGA��� ��{�CH�����TYPEm�y�a�[���� ��!JEW i������� �"////A/j/e/w/ �/�/�/�/�/�/�/?�?B?��WORD �?	p�
 	�RS��	�PNS2u��~2JO�
��TE[��?CO�Lu>8�?>L�� ��P��p���TR�ACECTL 1��Uz� .�`� ������|1LFDT Q��U�^@#@D � �sc/3BkO}I{O�O�D� �O�O�O�O�O_%__ _[]�Oe_�_9_�_�_ �_�_{_�^o�_�_To foxo*o<o�o@o�o�o �o�o
,>�i�a~�ccU� ����	���?� 1�S�e���i�����Ϗ �󏵏��+�=�O� �os�������џ��� ��+�=�O�a�s��� ��gI����ӯ���	� �-�?�Q�c�u����� ����Ͽ����)� ;�M�_�qσϕϧϹ� ��������%�7�I� [�m�ߑߣߵ����� �����!�3�E�W�i� {������������ ��/�A�S�e�w��� ������������ +=Oas��� �����'9 K]o����� ���/#/5/G/Y/ k/}/�/�/�/�/�/�/ �/??1?C?U?g?y? �?�?�?�?�?�?�?	O O-O?OQOcOuO�O�O �O�O�O�O�O__)_ ;_M___q_�_�_�_�_ �_�_�_oo%o7oIo [omoo�o�o�o�o�o �o�o�EWi {������� ��/�A�S�e�w��� ������я����� +�=�O�a�s������� ��͟ߟ���'�9� K�]�o���������ɯ ۯ����#�5�G�Y� k�}�������ſ׿� ����1�C�U�g�y� �ϝϯ���������	���-�?�Q�c��$P�GTRACELE�N  b�  ���a���w�_UP ��������В����w�_CFG ������a�
����������׉����DEFSPD� ���`щ���w�IN��TRL' �����8�F��PE_CONFI��Ш���t�����LID������	��LLB �1��� �t�B�  sB4��� ���� ���� 88�?�0�K�0� G�i�k�}��������� ����5Ak�����2���	�?��GRP� 1���lb�A�  �333a��A��D�@ �D�� D@ [A@�Ta�d+������� 	0='����´#��B 9!///O/�9/s/
��?�ö��/�/�.�/ =o=	7L�/ ?�/?P?;?t?_?�/��?�??�?�?�?  #DzC Oa�
OHO �?XO~OiO�O�O�O�O �O�O_�O_D_/_h_�S_�_�Z!a�
V�7.10beta�1�� Ax֝��R��y�Q?����Q>�\)f�QB0���PA��S�Bp���QA�9ASy�b
a�S �_`2oDoVoho��Ap���"���o�o�o�o����ө�KNOW_M�  ��֦�SV� ������5O8J\u_�@k}��Ҵ��M]��z�Д�R	��%%�"��|~���� ��u��P@�a�]�a�q�Xm��`��MR]��} ��&%O�P�$ӏ�K{ST]1 1���
 4��vi�Q:� �"�4�F�w�j�|��� ����ğ	����?�� 0�u�T�f��������P��ү��2� ��a��<K��^3 5�G�Y�k��4���������5ۿ���ς�6.�@�R�d��7 �ϓϥϷ��8�������
��MAD  �����OVL/D  ��G��PARNUM � ������T_S+CHy� ��
���8��0�UPD���������_CMP_0�p|�pp'�e��ER_CHK������j����RS8��oW_MO{����_���_RES_G��� o��� ������������ 2%VIzm`�R�4�\�l��Q���� ��S�ڰ�S� -�9X]S��x� �S������S�&���//S�V 1����a�q@c?\��THR_INRЮ�~��r�ed�&MA�SS�/ Z�'MN��/�#MON_QU?EUE ���fT"��a��N��U��qN�&��0END1;�79EXEF?75\��BEE0'?3OPT�IO$7D�0PROGRAM %�*�%0T/��2TA�SK_I{ԍ>OCFG ��/���?^"@DATA�s�+K��"�2��O�O �O�O�O�O�O_!_3_�E_�Oi_{_�_�_ROIWNFO�s�oM�
4 [_�_
oo.o@oRodo vo�o�o�o�o�o�o�o *<N`�W�T��oL �	!A�K�_%A�+I�^�vECNB|б})��v2���xG%A2��{ �P(O�4�F� �C�e��z_EDIT �+O����>DWERFLg8|#� �RGADJ M��:A����?"���!߆1�q�]�?�?���A<@��v%<�l�ӈ����q2�)��R	�H0le�{"6�?�
��AF$�t$�ܖ*�/� **:��"����� d�1�f�Ցd�[�_" U�#���3�E�s�i�{� ������߯կ�a�� �K�A�S�Ϳw����� ����9����#��+� ��O�aϏυϗ�߻� �������}�'�9�g� ]�o��ߓߥ������� U����?�5�G���k� }����-������ ����C�U���y��� ����������q -[Qc���� ��I�3);��_q���t&	 >O@/Հ./g/R$ݙ�/�ߓU/�/Q/�/�/�P?REF �)�Հ�Հ
߅IORI�TY�72F��MP�DSP�1яG7UT�FǓކODUCT�
A�:�/��OG��_TG΀B����2TOENT 1�� (!AF_INEq0OG?!tcpO6M�!ud%O^N!icmMOu��2kXY"�Í��X1�)� ��O�OX0��O�O�E�O)__M_ 4_F_�_j_�_�_�_�_ �_o�_%o7o*�3"���=Y�yo�o��>�+�J��/�io��o�������AK�,  �0�q'�9K]X5�7�pHA?NCE �)��rrn{d�o��uyw	3��?"3ق�POR_T_NUMr3X0����_CAR�TREPR0����SoKSTAq7 C��LGS @ȍ���K�X0Unothing�����̏�܌�����#��?k�T?EMP ɕ94�����_a_seiban�/���/�� ͟���ܟ� �9�$� ]�H�Z���~�����ۯ Ư����5� �Y�D� }�h�����ſ��¿�� ��
�C�.�g�R�w� �ψ��Ϭ�����	��� -��*�c�N߇�r߫� ���ߺ������)��M�8�q�\��6�k�VOERSIP0�7��� disab�le�r<�SAVE� ʕ:	26�00H844����,�!�.�@�_Od�C 	��{2 /����X�e����	-;
��c�n ��L��]_�0 1˧K�� "����0/URGE�pB�0T6l>5�WF� DOr6��r�6W�0�"�W�RUP_DELA�Y �;�R_?HOT %%&~1���+R_NORMALy�2���SEMI��"/�!_QSKIP���w�x��g/��/�/�/ r-�5�/�'�/??(? �/L?:?\?�?�?�?l? �?�?�? OO�?"OHO 6OlO~O�OVO�O�O�O �O�O_�O2_ _V_h_ z_@_�_�_�_�_�_�_����$RBTIF�?�RCVTMO�UT�B��`D�CR��E) ��~!B��D��5D!Z�A�F�� 6���r-�igĨ
��%���
�!�Ӆ�}/�o�f;�C�d;�pf<���<��.>�]�>П��o��o'8} 8^p ������� ���$�1%RDIO_TYPE  ��.�EFPOS1� 1���  x�����Ώ��� {����:�Տ7�p�� ��/���S�ܟ��� ՟6�!�Z���~���� =���دs����� ��� D�V���=�����¿ ]�濁�
ϥ��@�ۿ d�����#ϬϾ�Y�k� �����*���N���r� �oߨ�C���g��ߋ� �&������n�Y�� -��Q���u������ 4���X���|���)�;� u�����������B ��?x�7�[ �����>)b ��!�E��{ /�(/�L/^/�/ E/�/�/�/e/�/�/? �/?H?�/l??�?+? �?�?a?s?�?O�?2O �?VO�?zOOwO�OKO �OoO�O�O_._�O�O _v_a_�_5_�_Y_�_ }_�_o�_<o�_`o�_x�o�o|�2 1ш� 2oDo~o�o�o &oD �ohe�9�] ��
�����d� O���#���G�Џk�͏ ���*�ŏN��r�� �1�k�̟��🋟� ��8�ӟ5�n�	���-� ��Q�گu�����ӯ4� �X��|����;��� ֿq�����Ϲ�B�ݿ ��;Ϝχ���[��� �ߣ��>���b��� ��!ߪ�E�W�iߣ�� ��(���L���p��m� ��A���e������� �����l�W���+��� O���s�����2�� V��z'9s� ����@�= v�5�Y�} ���</'/`/��/ /�/C/�/�/y/?�/ &?�/J?�/�/	?C?�? �?�?c?�?�?O�?O FO�?jOO�O)O�O�o�d3 1ҵo_OqO �O)__M_SOq__�_ 0_�_�_f_�_�_o�_ 7o�_�_�_0o�o|o�o Po�oto�o�o�o3�o W�o{�:L^ �����A��e�  �b���6���Z��~� �����Ə �a�L���  ���D�͟h�ʟ��� '�K��o�
��.� h�ɯ�������5� Я2�k����*���N� ׿r�����п1��U� �y�ϝ�8Ϛ���n� �ϒ�߶�?������� 8ߙ߄߽�X���|�� ���;���_��߃�� ��B�T�f�����%� ��I���m��j���>� ��b����������� iT�(�L� p��/�S� w$6p��� �/�=/�:/s//��/2/�/V/�/�O�D4 1��O�/�/�/V? A?z?�/�?9?�?]?�? �?�?O�?@O�?dO�? O#O]O�O�O�O}O_ �O*_�O'_`_�O�__ �_C_�_g_y_�_�_&o oJo�_no	o�o-o�o �oco�o�o�o4�o �o�o-�y�M� q���0��T�� x����7�I�[����� ����>�ُb���_� ��3���W���{���� ��ß��^�I������ A�ʯe�ǯ ���$��� H��l���+�e�ƿ ��꿅�ϩ�2�Ϳ/� h�ό�'ϰ�K���o� �ϓ���.��R���v� ߚ�5ߗ���k��ߏ� ��<�������5�� ���U���y������ 8���\�������?� Q�c�������"��F ��jg�;�_����/45 1�?���n� ��f���%/� I/�m//�/,/>/P/ �/�/�/?�/3?�/W? �/T?�?(?�?L?�?p? �?�?�?�?�?SO>OwO O�O6O�OZO�O�O�O _�O=_�Oa_�O_ _ Z_�_�_�_z_o�_'o �_$o]o�_�oo�o@o �odovo�o�o#G �ok�*��` ����1���� *���v���J�ӏn��� ���-�ȏQ��u�� ��4�F�X����ޟ� ��;�֟_���\���0� ��T�ݯx�������� ��[�F�����>�ǿ b�Ŀ����!ϼ�E�� i���(�b��Ϯ��� ��ߦ�/���,�e� � ��$߭�H���l�~ߐ� ��+��O���s��� 2����h�������x9�16 1�< ����2����������� ����R��v �5�Yk}� <�`��� �U�y/�&/� ��/�/k/�/?/�/ c/�/�/�/"?�/F?�/ j??�?)?;?M?�?�? �?O�?0O�?TO�?QO �O%O�OIO�OmO�O�O �O�O�OP_;_t__�_ 3_�_W_�_�_�_o�_ :o�_^o�_ooWo�o �o�owo �o$�o! Z�o~�=�a s�� ��D��h� ���'���]�揁� 
���.�ɏۏ�'��� s���G�Пk������ *�şN��r����1� C�U����ۯ���8� ӯ\���Y���-���Q� ڿu�����������X� C�|�Ϡ�;���_��� �ϕ�߹�B���f�L�^�7 1�i��%� _�������%���I� ��F����>���b� �������E�0�i� ���(���L������� ��/��S��  L���l�� �O�s�2 �Vhz�/ /9/ �]/��//~/�/R/ �/v/�/�/#?�/�/�/ ?}?h?�?<?�?`?�? �?�?O�?CO�?gOO �O&O8OJO�O�O�O	_ �O-_�OQ_�ON_�_"_ �_F_�_j_�_�_�_�_ �_Mo8oqoo�o0o�o To�o�o�o�o7�o [�oT��� t��!���W�� {����:�Ï^�p��� ����A�܏e� ��� $�����Z��~���� +�Ɵ؟�$���p��� D�ͯh�񯌯�'�¯�K��o�
���yߋ�8 1ז�@�R���
� ��.�4�R��v��s� ��G���k��Ϗ�߳� �����r�]ߖ�1ߺ� U���y�����8��� \��߀��-�?�y��� �����"���F���C� |����;���_����� ������B-f� %�I��� ,�P��I� ��i��/�/ L/�p//�///�/S/ e/w/�/?�/6?�/Z? �/~??{?�?O?�?s? �?�? O�?�?�?OzO eO�O9O�O]O�O�O�O _�O@_�Od_�O�_#_ 5_G_�_�_�_o�_*o �_No�_Ko�oo�oCo �ogo�o�o�o�o�oJ 5n	�-�Q� ����4��X�� ��Q�����֏q��� ������T��x�����7�������MAS�K 1�û������XNO  ����MOTE�  3����i�_C�FG �p������PL_RANG�l�g�t�POWER� �õݠ|�S�M_DRYPRG %p�%m���TART �ծ�#�UME_PRO������_EXE�C_ENB  zd�x�GSPDX�우����TDB̽�ϺRM޿ϸI_�AIRPUR�� �p�B�<�ٛMT_��TРn��OB�OT_ISOLCB1��8�����9�z�NAME p��n�ۙOB_OR�D_NUM ?�ը5�H8�44 g���bҘ ����/(/�^/�Ҧ/���P�C_TIMEOU�T�� x�S23�2��1�4�γ �LTEACH PENDANP�X��������l��j�Mainte�nance CoKnsg��߾�"���f�No Use ���߮���0�B�T��h�NPO2�RҤ��z�e�CH�_L[��p���	����!UD1�:���R�VAIQL��R����x�e��PACE1 2�p�
 �濫��{鋓������9˺�?8�?�%��� %���4IDu� ������Y����� �):!4�8�Uu ������/ �):/!/O/q�� �U/���/ ?�/? 6??K?m//�/�/�/ c?�/�/�/�?O2O	O Oi?{?�?�?�?_O�? �?�OGO_._@_'_eO wO�O�O�O[_�O�O�_ o�_+_<o#oQos_�_ �_�_Wo�_�_�o�o 8Moo�o�o�o �o�o�o�D��4� �I�k}���a� ��돽��0�B��+�X�2a�s����� ��W�͏�����4�U�<�j�o�3~����� ��Ɵt����<��� Q�r�Y���o�4���� ��ѯ㯑��)�8�Y�@�nϏ�vϤ�o�5�� ʿܿ� Ϯ�$�F�U߀v�9ߋ߬ߓ���o�6 ����������A�c� r��V�������o�7����(�:���^� �����s���������o�8�!�3�E�W� {���������o�G �/� m�
u d  /��� ���/Nl -S -L/�/p�d� z ��/�/�/�/??&? /./@.1:n?�;�?�/ �/(?�?�?OO*O<O 2?D?V?h?�?�O�O�? �?HO__&_8_J_\_�ROdOvO�O�O�_ ` @p��U]/ o�O�IAakU�_Ro doj_DjEowo�o�o�o �o�o%�o�o= ASe���	� ��3�E���+�]����a�o\
#o�o�_MODE  /^
�S �/��_�Z�oH������	��㟐�CWOR�K_AD�
���D��R  /�< 1���_INT�VAL�a�%�R_OPTIONR�� %���V_D�ATA_GRP �2�uX:D�@P П��̟�˩͏��� 1��U�C�y�g����� ��ӿ������	�?� -�O�u�cϙχϽϫ� ���������;�)�_� M߃�qߧߕ߷����� ���%��I�7�Y�[� m����������� ���E�3�i�W���{� ������������/ SAwe�����P�$SAF_DO_PULS��Q�A��� CAN�_TIM��E}��R ���Ƙ�qsy�֡��Yo�K�C կ����� �l//%/7/I/[/Ve��C�2�$$K�)d�$�!ѢIf)�P5��/�/�/���)�/ ��4�w_ �R  T0��!?^?p?�?�9T D���?�?�?�?�?  OO$O6OHOZOlO~O �O�O�O�O�OU�s��'�O$_6_�I�  �T;��o��WQo�p�M
�?t��Di��[~=Z0 � �� o�[Q[SC�_�_�_ �_o o2oDoVohozo �o�o�o�o�o�o�o
 .@Rdv�� �������*��<�N�`�r�������� ?��я�����+� =�O���r%{������� ß՟�����"�_���02�SwU�]n��� ������ȯگ���� "�4�F�X�j�|����� ��Ŀֿ�����0� B�T�f�xϊϜϮ��� ��������,�>ߩ� b�t߆ߘߪ߼����� ���o�(�:�L�^�p� �����#�Q�[�� ��
��.�@�R�d�v� �������������� '9K]o�� ������# 5GYk}�������O�3�/ /1/C/U/g/y/�/�/ �/�/�/�/�/	??-?�;:�D?q?{6���d�j?@]	12345678�R�h!B!�U���B��V� �?�?OO)O;OMO_O qOwA��O�O�O�O�O �O__*_<_N_`_r_ �_�_�_�_�]�O�_ o o$o6oHoZolo~o�o �o�o�o�o�o�o�_ �_DVhz��� ����
��.�@� R�d�#��������Џ ����*�<�N�`� r���������y�ޟ� ��&�8�J�\�n��� ������ȯگ���� ϟ4�F�X�j�|����� ��Ŀֿ�����0� B�T�f�%��ϜϮ��� ��������,�>�P� b�t߆ߘߪ߼�{��� ����(�:�L�^�p� ����������� ����0.�@�%����l�~����Cz � B\�   ���2d4� ���d1
���  	�d22,�%X7IXp���Z������� %7I[m �������� !/3/E/W/i/{/�/�/ �/�/�/�/�/??/?@A?S?e?w?�?�:Z������<�4��`�$�SCR_GRP �1�� �� � ���� ��	 _�1��2 
BD[����� I�7GpDO2OkO������hBDE� DP��wC�GhK�A�RC Mate �120iC 67w890��M-�@�A 8��M2I�A�A��
123�45�D;F�2  ����>U�1{F�1 HC�1�AhAJ<ANY	?R�_�_�_�_�_~�\��H��0�T�7�2 o/O0oVoho7F/��Co�o?o��o���l0Q�o:DB�B���r2tAA���A  @��YuA@9�Wpj ?�wr�H��DzAF@ F�`�r��o� ����B�-�f�Q� ��}Yq�r������ďքB��y�*��N� 9�r�]�o�����̟�� �۟�&���CTOF�k�����h�����q�Yq>��̣�7G@hYpݯ����W \HC+�3���AnpC�HV��o~ec��W���� y���������pո��¿ P�(�%�7�I�v�b�SS���0EL_DEFAULT  m�_���u�?HOTSTR��d��u�MIPOWE?RFL  ����޶�WFDO�� ��� u�RVENT? 1���`��� L!DUM�_EIPL�(��j�!AF_INEx��Fߺ�!FTߒu�<ߙ�!o�� ������!RP?C_MAIN����q���1���VIS���ٻ �}�!TP&p�PUt�/�dl����!
PMON_POROXY��2�e�������+�f�a�!�RDM_SRV�b�/�gP���!R�T��0�h����!
���M,�,�i��E!RLSYNCF�l	84�!R3OS߸�4���!
CE��MTC�OM�2�k�)!=	�CONS*1��lu!�WA'SRC|�2�md�;!�USB�0��n�/!STM��'/.�o�Y/��}/ p�J/\/�/�/�/�/���ICE_KL ?�%� (%S?VCPRG1�/::"$52:???)03b?g?")04�?�?)05�?�?")06�?�?)07OO�)0
TJOE<9ROWK &4��O)1,?�O)1T? �O)1|?�O)1�?_)1 �?G_)1�?o_)1O�_ )1DO�_)1lO�_Q1�O oQ1�O7oQ1�O_oQ1 _�oQ15_�oQ1]_�o Q1�_�oQ1�_'Q1�_ OQ1�_wy1%o�/	2 )0?"0���1�/� �S�>�w�b������� я��������=�(� a�L�s���������ߟ ʟ��'�9�$�]�H� ��l�����ɯ��ۯ�� �#��G�2�k�V��� ����ſ���Կ����1��C�g�Rϋ��*_�DEV ���MC:��,����GRP 2��՟�0bx 	� 
 ,����ߟ���7��[� B�Tߑ�xߵߜ����� �����3�E�,�i�P� �������z������� ��A�S�:�w�^��� ������������+ O��D�<�� ����'9  ]D��z��� ��/h5/G/./k/ R/�/v/�/�/�/�/�/ ???C?*?g?y?`? �?�?�?�?*/�?�?O -OOQO8OuO�OnO�O �O�O�O�O_�O)__ M___F_�_�?x_�_p_ �_�_oo�_7oo[o moTo�oxo�o�o�o�o �o�oE�_i{ b������� ��A�S�:�w�^��� ����я�����^+� �O�a�H���l����� ��ߟƟ����9� � ]�D�����z������ �����5�G�.�k� R�������ſ����� ���C�*�<�yϟ�d ���	gϰϛ���Ͽ������+�%�x+�Pߌ����i� �i�y߇�qߧߕ��� ������=�"�e���O� =�s�a������� ��3��'��K�9�o� ]������������� ��#G5k��� ��[�W��� C�j�3�� �����/]B/ �/u/c/�/�/�/�/ �/�/5/?Y/�/M?;? q?_?�?�?�?�/�?�? �?�?�?OIO7OmO[O �O�?�O�?�O�O�O�O �O_E_3_i_�O�_�O Y_�_�_�_�_�_�_o Ao�_ho�_1o�o�o�o �o�o�o�oIooo@o sa����� !�E�9��I�o� ]��������ޏ��� ���5�#�E�k�Y��� я������ן��� 1��A�g�����͟W� �����ӯ	���-�o� T�f��?�������� �Ͽ�G�,�k���_� M�o�qσϹϧ���� �C���7�%�[�I�k� m�ߵ�����ߥ�� ��3�!�W�E�g���� ���ߍ��������/� �S���z���C���?� ��������+m�R ���s���� �E*i�]K �o����/ A�5/#/Y/G/}/k/ �/��/�/�/�/�/�/ 1??U?C?y?�/�?�/ i?�?�?�?�?�?-OO QO�?xO�?AO�O�O�O �O�O�O�O)_kOP_�O _�_q_�_�_�_�_�_ 1_W_(og_o[oIoo mo�o�o�o	o�o-o�o !�o1WE{i� �o������ -�S�A�w�����g� я�������)�O� ��v���?�����͟�� �ߟ�W�<�N��'� �o�����ɯ���/� �S�ݯG�5�W�Y�k� ����ſ��+���� �C�1�S�U�gϝ�߿ ��ύ������	�?� -�Oߥ��Ϝ���u��� ��������;�}�b� ��+��'������� ���U�:�y��m�[� �����������-� Q���E3iW�{ ���)� A/eS���� y�u�//=/+/ a/��/�Q/�/�/�/ �/�/??9?{/`?�/ )?�?�?�?�?�?�?�? OS?8Ow?OkOYO�O }O�O�O�OO?O_OO �OC_1_g_U_�_y_�_ �O�__�_	o�_o?o -ocoQo�o�_�o�_wo �o�o�o;)_ �o��oO���� ���7�y^��'� �������ُǏ��?� $�6����W���{� ����՟���;�ş/� �?�A�S���w���� ԯ������+��;� =�O���ǯ���u�߿ Ϳ��'��7ύ��� ��ÿ]Ϸϥ������� ��#�e�J߉��}�� �߳ߡ�������=�"� a���U�C�y�g��� �������9���-�� Q�?�u�c��������� �����)M; q����a�]� �%I�p� 9������� !/cH/�/{/i/�/ �/�/�/�/�/;/ ?_/ �/S?A?w?e?�?�?�? ?'?�?7?�?+OOOO =OsOaO�O�?�O�?�O �O�O_'__K_9_o_ �O�_�O__�_�_�_�_ �_#ooGo�_no�_7o �o�o�o�o�o�o�o aoF�oyg�� ���'���� �?�u�c�������� �#�����'�)�;� q�_���׏������� ݟ��#�%�7�m��� ��ӟ]�ǯ���ٯ� ���u���l���E��� ��ÿ���տ�M�2� q���e���uϛωϿ� ����%�
�I���=�+� a�O�qߗ߅߻����� !߫���9�'�]�K� m���ߺ��߃����� ���5�#�Y������ I�k�E��������� 1s�X��!�y� ����	K0o �cQ�u��� �#/G�;/)/_/ M/�/q/�/�/�// �/??7?%?[?I?? �/�?�/o?�?k?�?O �?3O!OWO�?~O�?GO �O�O�O�O�O_�O/_ qOV_�O_�_w_�_�_ �_�_�_oI_.om_�_ aoOo�oso�o�o�oo �o�o�o�o']K �o��o��� ���#�Y�G�}�� ���m�׏ŏ���� ��U���|���E��� ��ӟ������]��� T���-���u�����ϯ ���5��Y��M�߯ ]���q�����˿�� 1���%��I�7�Y�� mϣ����	ϓ����� !��E�3�U�{߽Ϣ� ��k����������� A��h�z�1�S�-�� ��������[�@������$SERV_MAIL  �����e�OUTP�UTt���RoV 2�	�  ��� (�O���i�S�AVE��g�TOP�10 2�� d ��;M_q ������� %7I[m� ������/!/ 3/E/W/i/{/�/�/�/ �/�/�/�/??/?	��YP��f�FZN_CFG �	�'��.��o1?GRP 2�y7��� ,B   A��0.D;� B��0�  B4.�RB21��HELLr2�	���������7"O1K%RSR1O2ODO}OhO�O �O�O�O�O�O�O_
_�C_._g_R_�_�_�^_�  ��%�_��_�_�R�\a. ��_b`ރ��R2�. do�_�6HK ;1��; o�o �o�o�o�o�o�o
3 .@R{v�������<OMM ���?2��2FTOV_ENBt�����HOW_REG_�UIR�g�IMIO/FWDL��!��5�A��*SYST�EM*. V8.3�0340 ł11�/9/2020 �A ���X��SNPX_ASG�_T   0 �$ADDRES�S  ��ZE��VAR_NAM�	�%$MULT�IPLY��P�ARAM�� � $TIME��v�$�_ID�	$NUM�D�T��CIMP[�FRI�FD�VERSIOyN��G�TATU ��$DISK�NF�OD�MODBUS�_ADR[�����P�ORC�`�SSR~�� x ���NGLE��g�$�DUMMY7�S�GL�TASK   &����T�x�����STMTT0��PSEGT2�B�WD�h��E��SVCNT_GP��� 8 $PC��ER_V�  � 	$FB�P�m�SPC��m�ΐV�DX�R[��� �$DATA0�Ӏ u���1��2���3��4��5��6���7��8��9��A*��B��C��D��2�B��F�� y���1ΩU1۩1�1��1�U1�1�1)�16�U1C�1P�1]�1j��1w�ҁJ���2Ω2�۩2�2��2�2��2�2)�26�2�C�2P�2]�2j�2�w�3��3��3Ω3�۩3�3��3�3��3�3)�36�3�C�3P�3]�3j�3�w�4��4��4Ω4�۩4�4��4�4��4�4)�46�4�C�4P�4]�4j�4�w�5��5��5Ω5�۩5�5��5�5��5�5)�56�5�C�5P�5]�5j�5�w�6��6��6Ω6�۩6�6��6�6��6�6)�66�6�C�6P�6]�6j�6�w�7��7��7Ω7�۩7�7��7�7��7�7)�76�7�C�7P�7]�7j�7�w���S�PRM�_UPDӑ � $4q� 
蛡��ӑؐ$T�ORQUE_CM�D   u�MO�a_SPEEjQ?_CURREo�nGAXI �mS��CART��_�Ut��̒YSLO~� � �@�����������_��{�VALU�OPб�$�#(F�ID�_L��K%HIF*I�N�$FILE1_A�v$�$M�t���SAR0  �h^� E_BLC�K���"���(D_CPU�)��)��F#y/�$���_=�R 	 � PWҐ�OT��)1LA#��SR� .3?184RUN_FLGQ5-4U184WITX5v1-4v1�85H2�D4�084|P��TBC2��
 O� $O�X0IG|u �0_FTM1D���42D�TDCX0A
Z��2M���6�1�7TH��C�DxG�R.0A��ERVE��3?D�3?D3O��0_�AC@ Xw -$jALEN�3�wD�3j@EL_RA�TI��$�W_��F#1jAc$2�GM�O�!>��C��ERTIA�o!�Iaj@�K�DE�E��LACEMM�CC�CmV�@�MA��F7UW7QT�CV>\_QWTRQ ^\UuZ���Ct��US&t�J_��q�M�TF��J2'���E�QUvA2�P>�s�a�C@JKfVK�1'a�1�'a`A`J0<d+cJ�J3cJJ;cAAL�+ca`3ca`[f4\e5C�PN1�\�`Q[;PJ�L�@_�E��3�CF� `^G�ROU1 ����y�N��0CC��`REQUsIR*B��EBUZ��fA�V$T�@2�#qg@v�14 }\�ENABL	��$APPRpC�L�
$OPEN�`xCLOSEozS�E�y�E
�1.� �u M�0<PPB�t'_MGr!�pC��� p�x��9P�wBRK�y�NOLD�vh�RT�MO_�3���uJ"��PcdP3cP;c PcP�cP6P��S�b� @@eB�4�� r�B�1x���1��PATH���ӁɃӁ�Hσ0�(p�W�SCATr�ar6�qINiBUC�@��Z)�C��UM2�Y�@+@�P9�O!EAT��0�T�`@T�PAYLO�A�J2L7R_AN�1��L*0����������uR_F2LgSHR9DؑLO���(�ٗF��F�ACRL_�!&��"���B9H$ �$H�rG��FLEXcs�1J�6 PMr�?�?>O�PO�"d�iE :vO�FP٧�OA0P�O�O�LF1�>� R��O�O�O�O_!_��E+_=_O_a_s_�_�_ �_�_Y�vĽW�Sdf�@���_�_ o�jT2'W�X�`�eŴ��e '� �*o<oNo``deme [ee�o�o�o�i/d��d ��0�o�o�� 8ATk�q�PE�Lٰ}1=�xJ(pv#pJE �CTR"��f�TNR9�wHA_ND_VB�c��0 �� $��F24�v	D#SW�"�2��v� $$M ���yv�q���q�����>��AR ���vQ!D5��}A�| �zA�{AA�@��{� �zD�{�D�P�G@0��S�T�w���y��N�DYW0^p�v!�H���k@ ϗ�ϗꑎ�g������PX�a�j�s�|���������ӵ5 ���Ť����qA'SYM��^�p��!����_�0� .�A�+�-��K�]�o�����J��K�����\˙x�_VI��	(|�s V_UNIC.$P�בJeG"uG" �K$�X$|&
��P� K�,�>��%�T�\���1�0H+0Rr0���!v�VrDI�s�O4��� �c `�O�I2AO�F�I1 l�WW3o��1�۱�   � ��ME��@r2�"YT0PT���ڀ�1�`��u���8�1�9�T��a $D�UMMY1`A$7PS_i�RF+����$�6XpFLA��`YP��B�3$GLB_T��5*E��0Vq�`��j�v1 �XMpw��ST±�#pSBR��M21�_VrT$SV_�ER��O� pC�CC)LD@pBAڰOL2� �GL EW� �4�`�1$Y��ZB��W�C`ԑ��As0�2��"�@U�E ���N�@�$G�Iz�}$�A p�@�C�@� L�`\V�}$F�EV�NEAR��Np�F<]Y��TANCp��!�JOG�A� ���$JOINTx
����EMSET�  WECU۱��S���*R��׼ g�U��?��#pLOCK_FOx���0BGLVm��GLhTEST_sXMcp�QEMP�P�r+bBB�P$U���B2�2#p�CQa�b���PQarAC�E�`Sr` $KA�R�M3TPDRqA�@�d�QVEC���f�PIUQaVaH=E�PTOOL2��c�V1�RE�`IS3䱥�b6s�f�ACH�P(p�aO��3�4�29�2�`ISr � @$RAIL_�BOXE
��@R�OBO"d?��AHOWWARO�Aq�0qROLM�2gu���
txr��/pZ���O_=F��! �D�a�� �_ �R�`OBˢ!�r*��Q�p�FKOU�R"XBMeY�C���P$PIP#fN���b/r�ax�Qa��p��CORDED��P��q� ��OY0 �# D )@OBu�G��Pd�S��3(@�S��I�SYSS�A�DRH�� �0TCHl�S� ,0EN2*�A�Q_T���Ѽ��� VWVAu1% � �`�B5PREV_RT��$EDIT�V/SHWR��\F$�����A	 D�0���;���$HEADД� U���KE|�A�0CPSPDl��JMPp�L5b�R���44&[�t���Ij,`SH�C��NE�`<I��TICK2�<eM}��!��HNRA' @]�����t��_GP�&v��STY��qLODA�C��|��m�( t 
 �MGƅ%$�T=\@S>�!$=!2��1�EF0FP�SQ�U�`%�B!TER�C�0��TS��) Ph@�׹��׈g��a�`O�0�3t�I�ZDQE�1PR`E��1!����pPU��1�_DObR��XS:�PK6AXIP��sVaUR�ڳI�Hp��~����_�`��EET��P bl�O��FP�A��4 ss`��BSR��*lѠ��A� �������#�� 1��A�R�c�R�s�R� ��d�~Ͱ�dŢ������ː�C��|����SC,@ + h�@DS��a�03SPC0~�ATq���2�𐿒�2ADD�RES�cB�SH�IF�H`_2CH�H�z�IK@���TV�I72,��h��T�� 
+j
��V�q�A���- \���� O����<�C���൲���B<��TX_SCREEU�.	0=k�TINA�CP���T�A����� / T���@����Ag@���^���^����RROL wP��f���v��A;UE��0 �� ��r@S�A��RSM�T�UNEX��6F�� S_�Cf�6V�i����6��C�RB��� �2/��UE�1p=2�B��!�GMT� �Li!m�w@O�WB�BL_pW�0��2S �O�O�AcLE��GpTO�3�RIGH&BRyD�D��CKGR�0�NTEX��OJWIDTHs1�u��1�A�a%�I_�0H>�� 3 8�!wP!_T��ҭ�0R�@�R sw�2$� O�ѭ�%4���GG U2 �9R brqLUM�u����ERV
��@� P�aP�У5{0�G�EUR&cF���Q)&]�LPM��E��C�)jS�x�x�`wU5u6u7u8Z����3�9P��6�a��QS��4�US=R�D6 <���0qUR��RFOC�a.PPRIαmp�!�L TRIP+qm��UN$0547	P t�$0��Yq��Hb����� 8�  �G �\�T�p1��ѣ"O	S�1�&R���#�a�9�O�C�N�"�$�IaUU�:�/�/�8U��#OFF!`���;[�3On0 �ٰW5�4:�@GU�Nw��0B_S�UB�2p@��SRT�� �<��vQ�p �O9Rp�5RAU��4�T�9���1_���=s |���OWN� >T$SRC����r�D!`CE�MPFqI*�*ё�ESP-� �����e*B�&�b�!�B���> `10W�O8�T�COMP:1$��� _^@��b�A�q�EWA�C�?a�A�@�C�A�C ��VCCH�? ��qC36MFB1����qVC4�Y`��@�x %rT��� XdP^��spC�pRU�DRIV���_�V�uT̐fpD�MY_UBY�ZTV�񕠧�B��X�a�RGP_Sp�+��RL7��BM$��DE�Y��EX����EM�U��X7d[�US�P�po��<1G��P�ACINΑ}�RG MAadwbF3wb3wb���ARE����a�rH6Twb�pA R�@G�P�Pr�a6UR� �pBC d�_���2	�B�N�RECcSWo`_IApa�8c�O!���A��1s�E�U�B�� �q$7THKG�C��Iz���.p��zsEA���w�@x� 1u5UMRCV��WD �FOS�M� �Cs�	�rX3�c�rREF���v�v�q p7 ��p �z��z��{;��vp_@@�zq��{��S�/g�S�6�8R��E �$�=�ߠ4) �UӠOU��b<�ZS @�e2х2�$��R� �ΐ�B��2Ѻ�Kq�SUmLs�C�@CO:�f� D)`�NT�C Z��BY��e�!e�$�L�S���S�����!��JTǤFt �+��ǱT� ��CACH+�LO�����*`����@ܣC_L�IMI��FR%�T8j�'���$HO� 6B=�COMMpSB�O0 ]�Ԉ�I؄h@�VP�b����_SZ�3n���6����12 ���[`��&����Aa�MP�FAI&�G�vt��AD��BM�REׄ9�_SIZ��PH�`��FAS�YNBUF�FVR�TDk�w�I�aOL���D_@3��W3PN�ETUc�QNp�[�ECCU�hVE�M�`��۲&�VIR9C���VTP�pO���J�s�A�w�_DEcLA�cP�ƪŕ���G�p9pCKL+AS�3	ő_�F��ƀHp"�S;��N���PLEXEEI���B/��3cFLK I `]�^A��M��Ȅdws�.�^@�bJ# �ʱ��#�#RS. ORD@!��> �3 ނ)�K��TB\"���WwCb2V��g%L`�Qۑ6D4���\*bUR3cp_R '�d���,a]��ծc�_ od&�{g��`B*�9T�'�SCO��*�C� ad�"_f�"0�" >�"K�"Y�J_\_nZh��� E\ AM�Pn�0 PSMf%sMp"%HADJT�F/e��Bڒ� Np"�q׬!LIN]3q���XVRh$O\���T�_OVR� �ZABC�5P�bw�$Ӻ�
O�ZIPg%Q�p"DBGLV�CL��R ���MPCF��5R  r ���$\��QLNK�2
��-`|�S �|q�����CMCMi`C�CC��ACtP_�  O$J:4D�� @QJ�V�4$08�tO�UXW� ��UXE>a��E��[���	���=Z��T ���Ԫr�YK�D"0 �U�"��^IGH�bcq�?( �K��|V � vG��$B$��@1e�B��,��&GRV%�F� ���OVC�5�A7�Pw@�`��
VBI����D�TRACE�B�V;1SPHE}R�P W , ��3I[�$SIM��A-Q��e!4P �`e!V&��qe!�m/!��%���/Kpb/�t#_UN�@_+�p&LCд�% ��%V M��ALI�AS ?e����%1�! ( he�!:?L?^?p?�?�6 6?�?�?�?�?�?	OO -O?OQO�?uO�O�O�O �OhO�O�O__)_�O M___q_�_._�_�_�_ �_�_�_o%o7oIo[o oo�o�o�o�oro�o �o!3�oWi{ �8������ �/�A�S�e������ ����я|�����+� ֏<�a�s�����B��� ͟ߟ����'�9�K� ]�o��������ɯۯ �����#�5��Y�k� }�����L�ſ׿��� ϸ�1�C�U�g�y�$� �ϯ�����~���	�� -�?���c�u߇ߙ߫� V�����������;� M�_�q��.����� �����%�7�I��� m��������`����� ��!��EWi{ &������ /AS�w�� ��j��//+/ �O/a/s/�/0/�/�/ �/�/�/�/?'?9?K?�]?3�$SMON�_DEFPRO �����1� *S�YSTEM*p:R�ECALL ?}��9 ( �}�tpdisc 0�=>172.8.�9.225:13�524 4  m�d: over �=>351928�32:10268�8d?O"O2L}t�pconn 0  �?�?�?�O�O�O;G�? WOiO{O__0_�BHB1�O�O�O�_�_�_�O �O^_p_oo%o8OJO��_�_o�o�o6l9c�opy virt�:\output�\untitle�d1.pcdovb6�975�o"5m7��bfrs:ord�erfil.da�t�dtmpback\�_4 �o���4n.�bmdb:*.*[Qnu��*�6=e2xFt:\�P��4 �������Aa3F�aN�`��u{����0� }
xyz�rate 11 �я���������=e<F�f�7864P�f� x�	��-�@b�_ږ �󟄯����;oMl\� n����#���:�o�o�jc1917583�36:16538!62�������6FXBN� }�� ϳ�-���ٗ���ϗϩϼ�1 F�Y�՛x�	��-�@� Ώ��ܔ�ϊߜ߮�A� S�e�w���,�?��߀���߆��｟M\4092 c�u��� *�=������������ ��Ml\�n���#6� H��������������968bt)<�� ���� �����]o //$/ 7I����/�/��Wb�`6b/t/??)?<�/ �/�/�?�? �?�Ml\?n?�?O#O����Z��28802�2784:9515802O�O�O��ȿ ڿ�.}O_ _�OE��O �(�O�_�_�_��O�a� �#x_	oo-o@��_�_ � �_�o�o�o�O�O\_ w_,?_Q_c_�o����;D�$SN�PX_ASG` �����q�� P 0 '�%R[1]@g1.1��y?�;C%�(��L�/�A��� e�������܏��я� ���H�+�l�O�a��� ����؟����ߟ�2� �<�h�K���o���¯ ��̯��ۯ����R� 5�\���k�������� ſ����<��1�r� U�|Ϩϋ��ϯ���� ���8��\�?�Qߒ� uߜ��߫�������"� �,�X�;�|�_�q�� �����������B� %�L�x�[�������� ������,!b El�{���� ��(L/A� e������/ �/H/+/l/O/a/�/ �/�/�/�/�/�/�/2? ?<?h?K?�?o?�?�? �?�?�?�?O�?ORO 5O\O�OkO�O�O�O�O �O�O_�O<__1_r_ U_|_�_�_�_�_�_o �_o8oo\o?oQo�o�uo�o�o�d�tPAR�AM �u��q �	��jP�;tAp�h#t���pOFT_KB_?CFG  s�u��sOPIN_SI/M  �{vu���p�pRVQS�TP_DSB^~�r��x�`SR �ay � & SOCKET��"��vTOP_�ON_ERR  �-�Kx?�PTN ��fr�A�;�RING_PR�MI� �`VCNT_GP 2au:&q�(px 	�̏�p���ޏ��wVD>��RP 1�i'p�y�R�d�v��� ������П����� *�<�N�`��������� ��̯ޯ���&�M� J�\�n���������ȿ ڿ���"�4�F�X� j�|ώϠϲ������� ����0�B�T�f�x� �ߜ߮���������� �,�>�e�b�t��� ����������+�(� :�L�^�p��������� ������ $6H Zl~����� �� 2DV} z������� 
//C/@/R/d/v/�/ �/�/�/�/�/	??? *?<?N?`?r?�?�?�? �?�?�?�?OO&O0��PRG_COUN��At�r�NuRBENB��MEMwCAt�O_UPD 1�{T  
;Or�O �O�O__(_:_c_^_ p_�_�_�_�_�_�_�_  oo;o6oHoZo�o~o �o�o�o�o�o�o  2[Vhz�� �����
�3�.� @�R�{�v�����Ï�� Џ����*�S�N� `�r����������ޟ ��+�&�8�J�s�n� ��������ȯگ��� �"�K�F�X�j����� ����ۿֿ���#���0�B�k�f�x�DL_I�NFO 1�E��@��	 �����������@��@�@�>�����.�
� �������A�/���%q���w�Av����o߁� Da���q~D��Q�6���´��ߞ�O@YSDEBSUG\@�@��d�I���SP_PASS�\EB?��LOGW ���C��9�ؘ�  ��A��UD1:\�<���_MPC�EH���AH�� �A~m�SAV �m�4�L��S�S�Vd�TEM_TI_ME 1	��@W 0����Ā���_��$T1SVGgUNS�@]E'�E��r�ASK_OPTION\@�E�A�A��_DI��xO���BC2_GRP �2
�I=�����@��  C�f�BC?CFG ����s l�]`] `ߕ������ �7"[FX� |������/ 3//W/B/{/f/�/�/�/�/���,�/�/"? 4?�/?j?U?�?y?�? ���?���0�? O�?$O OHO6OlOZO|O~O�O �O�O�O�O_�O2_ _ B_h_V_�_z_�_�_�_ �_�_�_�_.oh� Bo Toro�o�oo�o�o�o �o�o&8\J �n������ �"��F�4�j�X�z� ����ď���֏��� ��0�f�T���@o�� ��ҟ���t���*� P�>�t�����f����� �ί����(�^� L���p�����ʿ��ڿ  ��$��H�6�l�Z� |�~ϐ��ϴ��Ϡ�� �2�D�V���z�hߊ� �ߞ����������
� @�.�d�R�t�v��� ���������*��:� `�N���r��������� ������&J �b t���4��� �4FX&|j �������/ /B/0/f/T/�/x/�/ �/�/�/�/?�/,?? <?>?P?�?t?�?`�? �?�?OO�?:O(OJO pO^O�O�O�O�O�O�O  _�O$__4_6_H_~_ l_�_�_�_�_�_�_�_  ooDo2ohoVo�ozo �o�o�o�o�o
�?" 4Rdv�o��� ������<�*� `�N���r�������ޏ ̏���&��J�8�Z� ��n�����ȟ���ڟ �����F�4�j� �� ����į֯T����
��0��T�>�r��$T�BCSG_GRP� 2>���  �r� 
? ?�  ���� ��ӿ������-���Q�c�v�}���d�0 ���?r�	 HC�`�r���~b�C�  B�x���Ȣ�>�ff��"�ƞ�������϶�e\��H �h�BLc���B$дh�j߈� �߲߰����ތ��@�@��AƷ�f�y�D�V�������	��?�333��2�	�V3.00��	�m2ia�	*�T�L�q�c�"���e�r����� ��|l���   ��aB������u�J2}����5���CFG� >��� ,��
�D��Go�o��
G� ������5  YDV�z�� ����/1//U/ @/y/d/�/�/�/�/�/ �/�/????Q?���� \?n?�?*?�?�?�?�? �?O�?1OOUOgOyO �OFO�O�O�O�O�O	_ r�^�._:�>_@_R_�_ v_�_�_�_�_�_�_o *ooNo<oro`o�o�o �o�o�o�o�o8 &\Jl���� �������6�X� F�|�j�����ď��ԏ ����܏.�0�B�x� f�������ҟ����� ��*�,�>�t�b��� �������ί��� :�(�^�L���p����� ��ܿʿ ��$��H� 6�X�~�(��ϨϺ�d� ���������D�2�h� Vߌߞ߰��߀����� 
����@�R�d��t� ������������ ��*�`�N���r��� ����������& J8n\~��� ���"��:L 
�|���� ���0/B/T//d/ �/x/�/�/�/�/�/? �/,??P?>?`?�?t? �?�?�?�?�?�?OO OLO:OpO^O�O�O�O �O�O�O�O_ _6_$_ Z_H_j_l_~_�_.�_ �_�_�_ oo0oVoDo zoho�o�o�o�o�o�o �o
@.Pv� �Tf����� �<�*�L�r�`����� ����ޏ̏����8� &�\�J���n������� ڟȟ���"��F�X� op���o>�į��� ֯����B�0�f�x� ��H�Z������ҿ� �,�>���b�P�r�t� �ϼϪ��������(� �8�^�L߂�pߦߔ� �߸�������$��H� 6�l�Z��~����� ��d����&�����D� V���z����������� 
.��R@bd v������ *N<^`r� �����//$/ J/8/n/\/�/�/�/�/ �/�/�/?�/4?"?X? F?|?�?8��?�?�?t? �?�?OO.O0OBOxO fO�O�O�O�O�O�O�Op__>_(^  dP�hS hV|_hR��$TBJOP_G�RP 20U��  ?��hV	�R�S�\��8P���p��Q�U  � � � ��R�hS @dP�R	� �C� ff�  C�W�Q4b�<f9o >�f�f\a<a=�ZC]�`���b�&`�H&`.g�o�gn�`�W4e\e`b�o ?a~�d=�7LC�no#BȂo#&`�`9u�o�c�33\uX2h~�P<��C\vc�@333@330|b}`�BL�wHqsDa�l����u��Jh�p<X��B�$�d��?���C*p��C����Z`y�x��k< ���q`?]`C4�.�ϏR�d��daG�x���{<g����]p@&b`yap� c�z{4ep�V����� �����ʟ���(��  �N��Z��������P��ޯ��d�hV0��4e	V3.00��Sm2ia�T�*Z��TcQh�s� �E�'E�i��FV#F"w�qF>��FZ�� Fv�RF�~�MF���F����F��=F����F�ъF���3F���F��{G
G�dG�G#�
��D��E�'
EMKE����E�ɑE��ۘE��E����F��F���F��F(���F5��FB���FO��F\���Fi��Fv���F��vF��u�<#�
<Kt���@Ť�r_X�j�M�hTn�@�U��S��SESTPARaSA�\X�P�SHR��ABLE 1�[I��hS�ȃ� �0cɞ�����gWoQ*��	��
������*hQ������C�N��RDI�ϬQ��@� �2�D�Vվ�O�߀��������*���S�ߪS �������!� 3�E�W�i�{������� ��������/A �]�����̂	k�}�� ��M�_�q߃ߕߧ���~hNUM  0U��Q�PpP �B�C���_CFG �P�a@�PIM?EBF_TT���8�S���VERAÔz��R 1�[O 8e�hRcP2! 3P�  � / /$/6/H/Z/l/~/�/ �/�/�/�/�/�/? ? 2?{?V?h?�?�?�?�?��?�?�>��?O�: 0OBOTO.OxO�OdO�O �O�O�O�O�O_,__P_b_�8�_�_�_~_@�_�_�_�_���_K��@���MI_�CHAN� � >mcDBGLV逡����p`ETHE�RAD ?��
�`�n��?o�o�o���p`ROUT��!p
!"t@|SNMASK�h��a255.~uF�|���F���OOLO�FS_DI��GT ��iORQCTROL p	��n��T�B�T�f�x��� ������ҏ����� ,�>�P�b�r�����������PE_DET�AI�h�zPGL_�CONFIG �Qa��/c�ell/$CID?$/grp1��3� E�W�i�{�1�	�� ��ʯܯ� ���$�6� H�Z�l�~������ƿ ؿ�������2�D�V� h�zό�ϰ������� ��
ߙ�.�@�R�d�v� ���)߾���������}��N�`�r��@�������턬� ��)�;�M�_��߃� ����������l� %7I[m���� ����z!3 EWi����� ����///A/S/ e/w//�/�/�/�/�/ �/�/?+?=?O?a?s? �??�?�?�?�?�?O �?'O9OKO]OoO�OO �O�O�O�O�O�O_���User �View !�}}�1234567890B_T_f_x_�_�_��T-`��_��(Y2 5Y�Ooo*o<oNo`o�_�_/R3�_�o�o�o@�o�ogo)�^4�o bt������^5Q�(�:�L�^�p�����^6�ʏ܏�� ��$���E��^7 ��~�������Ɵ؟7����^8m�2�D�V�h��z���럭��� �lCamera3Z)����(�:�L�*�E�v�����@_���ƿؿ�����  ̦�Y�^�pςϔ� �ϸ�_����� �K�$�@6�H�Z�l�~ߥ��̦ �i������� ��$� ��H�Z�l�ߐ��� ������ߣ�Py��6� H�Z�l�~���7���� ��#��� 2DV ���*������� ����"4F�j |����kͥ�� Y/ /2/D/V/h/ �/�/�/��/�/�/
? ?.?���l��/z?�? �?�?�?�?{/�?
OO g?@OROdOvO�O�OA? �� �1O�O�O
__._ @_�?d_v_�_�O�_�_@�_�_�_o�O�G9�_ GoYoko}o�o�oH_�o �o�o�_�o1CU(gy�	Υ0�o� ������o2�D� V��oz�������ԏ {�Ӡիx�-�?�Q� c�u���.�����ϟ� ���)�;�M��Υ A�䟙�����ϯ�� ���)�;���_�q��� ������`��u��P�� �)�;�M�_���ϕ� �����������%� ̿޵���q߃ߕߧ� ����r�����^�7� I�[�m���8�޵� (�������%�7��� [�m����������� ������޵���I[ m��J���� 6!3EWi  	��� ���//(/:/L/^+   nv�/ �/�/�/�/�/ ??$? 6?H?Z?l?~?�?�?�? �?�?�?�?O O2ODO VOhOzO�O�O�O�O�O �O�O
__._@_R_d_�v_�_�_�_�_�_b, � 
 (  �>�( 	 �_o o:o(o^oLo�opo�o �o�o�o�o �o$�Z~* ̸i{ � ������ X5�G�Y��}��� ����ŏ׏����� f�C�U�g�y������ ��ӟ�,�	��-�?� Q�c������������ ����)�;���_� q���ʯ����˿ݿ� �H�%�7�Iϐ�m�� �ϣϵ���� ���� !�h�E�W�i�{ߍߟ� ��������.���/� A�S�e�߉����� ��������+�r�� a�s������������ ��J�'9K��o ������� X5GYk}� �����0// 1/C/U/g/��/�/�/ ��/�/�/	??-?t/ Q?c?u?�/�?�?�?�?p�?�?:?p@ B�"O4OFOCG `���)frh:\t�pgl\robo�ts\m20ia�\arc_mat�e_1�@c.xmlO�O�O�O�O�O_`_(_:_L_XX��X_ }_�_�_�_�_�_�_�_ oo1oCoZ_Toyo�o �o�o�o�o�o�o	 -?VoPu��� ������)�;� RL�q���������ˏ ݏ���%�7�N�H� m��������ǟٟ� ���!�3�J�D�i�{� ������ïկ���� �/�F�@�e�w����� ����ѿ�����+�t=�_H�1 O�j@88�?� =�|�=�xϚϜϮ��� �����0��<�f�P� rߜ߆ߨ��߼�����&��$TPGL_�OUTPUT �"H1H1 `�H�]�o���� �����������#�5� G�Y�k�}����������������H�`���2�345678901 2DVhz� >2����� �9K]o�}������� �1/C/U/g/y/�/#/ �/�/�/�/�/	?�/? ??Q?c?u?�??1?�? �?�?�?OO�?%OMO _OqO�O�O-O�O�O�O �O__�O�OI_[_m_ _�_�_;_�_�_�_�_ o!o�_/oWoio{o�o �o7oIo�o�o�o /�o=ew��� E�����+�� �}[�a�s����������̍@b����h�? ( 	 7� %�[�I��m������� ��ǟ���!��E�3� i�W�y�����ï��� կ�����/�e�S����^�w���ѽ �����)�;��� d�v�ϚϬϊ����� L���ߺ�(�N�,�>� �ߖ� ߺ���n���� ��&�8��D�n��^� ��������V��"� ��F�X�6�|�����z� ����x�����0B ��fx���� �N`,�Pb @����p� /�/:/��p/�/ $/�/�/�/�/�/X/�/ $?�/4?Z?8?J?�?�? ?�?�?z?�?O�?2O DO�?POzOOjO�O�O �O�O�ObO_._�OR_ d_B_�_�__�_�_�_��_oo�_<oNoTb��$TPOFF_L�IM ���p�����qibN_S]Vm`  ӄj�P_MON #����d�p�p2�ӅiaSTRTCHOK $��f^���bVTCOMPA�T�hq�fVWVA/R %�mAx�d� �o Y�p��bia_DEFP�ROG 3vb%?SOCKEp���m_DISPLA�Yt`�n�rINST�_MSK  �|� �zINUSE9R�tLCK��{�QUICKMEN�A��tSCRE`����rtps�c�t�{���b��_敉STziRAC�E_CFG &��iAtx`	bt
�?�܈HNL 2E'�i}� �H{ nr 4�F�X�j�|��������ĚޅITEM 2�( � �%$1�23456789y0��  =<�x7�I�Q�  !W�_�kp���bs�ů )����_������^� ��y�ݯ����5�%�7� I�c�m�翑�=�c�u� ٿ�����!ϛ�E��� �)ߍ�5߱�����Y� �������A���e�w� @��[�����ߧ� �k���O��s��E� W���c������}�'� ����o�/������ ;S����#�G Y"}=�as� ���1�U/ '/������_/ 	/�/�/�/Q/?u/�/ �/?�/i?�?�??�? )?;?M?�?O�?COUO �?aO�?�?�OO�O7O �O	_mO_�O�Ol_�O �_�O�_�_�_3_�_W_ i_{_�_�_Koqo�o�_ �ooo/o�o�oeo% 7�oC�o�o��o� ��O�s�N��ڄS�)�S��g  ϒS� �����y
 ��ݏď����UD1:\����e�R_GR�P 1*��� 	 @�pY�k��U���y�����ӟ��� ����͑�2��V�A�?�  q���m� ����ǯ���ٯ���� �E�3�i�W���{��������	!����~c�SCB 2+o� \�Y�k�}Ϗ���ϳ�������Y�V_�CONFIG �,o�󁧏�M���O�UTPUT -<o�>���Yߝ� ����������	��-� ?�Q�c�u�;ъߝ�� ��������	��-�?� Q�c�u���������� ����);M_ q�������� %7I[m �������/ !/3/E/W/i/{/��/ �/�/�/�/�/??/? A?S?e?w?�/�?�?�? �?�?�?OO+O=OOO aOsO�O�?�O�O�O�O �O__'_9_K_]_o_ �_�O�_�_�_�_�_�_ o#o5oGoYoko}o�_ �o�o�o�o�o�o 1CUgy�'�9� �������#�5� G�Y�k�}������oŏ ׏�����1�C�U� g�y���������ӟ� ��	��-�?�Q�c�u� ��������ϯ��� �)�;�M�_�q����� ����˿ݿ���%� 7�I�[�m�ϑϣϴ� ���������!�3�E� W�i�{ߍߟ߱����� ������/�A�S�e� w����������� ��+�=�O�a�s��� ������������ '9K]o��� ������#5 GYk}����x������ �/�3/E/W/i/{/ �/�/�/�/�/�/�/? �/?A?S?e?w?�?�? �?�?�?�?�?OO*? =OOOaOsO�O�O�O�O �O�O�O__&O9_K_ ]_o_�_�_�_�_�_�_ �_�_o"_5oGoYoko }o�o�o�o�o�o�o�o 0oCUgy� ������	�� ,?�Q�c�u������� ��Ϗ����(�;� M�_�q���������˟ ݟ���%�6�I�[� m��������ǯٯ� ���!�2�E�W�i�{� ������ÿտ������,��$TX_S�CREEN 1.����}ipnl/`�gen.htm,��ϑϣϵ���$ �Panel se7tup��}���� �0�B�T�f����� �߯���������n�� ��?�Q�c�u���� "���������)��� ����q����������� B���f�%7I[ m��������� �t��EWi{ ���:��/�///A/�/�UAL�RM_MSG ?5L��Y� Z//� �/�/�/�/�/�/?? $?B?H?y?l?�?�?�?~u%SEV  �-��6s"ECFG� 0L�V� � /�@�  A�#A   B�/�
 �?6�L�VOhOzO �O�O�O�O�O�O�O
_�W�1GRP 21�	K 0/�	 �@Ob_u I_BBL�_NOTE 2�	JT���l6�Q�8�@uRD_EFPRO %�+ (%�?�_8��_ o�_'ooKo6oooZo��o�o�o�o�o�ok\I�NUSER  ��]P_�oI_MENHIST 13	I  ( �P���(/SOFT�PART/GEN�LINK?cur�rent=men�upage,153,17����<o�,195�,��>�P�b��p'��7�1�����ӏ��q+�y��edit�rSOCKET��7�I�0[��x���34&��� ɟ۟��q�o�'�9� K�]�o���������ɯ ۯ�|��#�5�G�Y� k�}��Rlq�����Ϳ ߿���'�9�K�]� oρ�ϥϷ������� �ώϠ�5�G�Y�k�}� ��߳���������� ��1�C�U�g�y��� ,���������	���� ?�Q�c�u��������� ������),�M _q���6�� �%7�[m ���D��� /!/3/�W/i/{/�/ �/�/�/R/�/�/?? /?A?�/e?w?�?�?�? �?�����?OO+O=O OOR?sO�O�O�O�O�O \O�O__'_9_K_]_ �O�_�_�_�_�_�_j_ �_o#o5oGoYo�_}o �o�o�o�o�o�oxo 1CUg�o�� �����?�?�-� ?�Q�c�u�x������ Ϗ�󏂏��)�;�M� _�q��������˟ݟ ����%�7�I�[�m� �� ���ǯٯ��� ���3�E�W�i�{��� ���ÿտ��������$UI_PA�NEDATA 1�5���A��  	�}�/frh/cg�tp/wided?ev.stm�z���Ϟϰ���)prih��ϧ�}���"�04�F�X�j� )lߐ� wߴߛ���������� 2�D�+�h�O�������� �  ��M� �����#�5�G�Y��� }��ϡ����������� b�1U<y� r�����	� -?&c�� D�� CÞ������� P!/��E/W/i/{/�/ �//�/�/�/�/�/? /??S?:?w?^?�?�? �?�?�?�?Oz�=O OOaOsO�O�O�?�O./ �O�O__'_9_K_�O o_V_�_z_�_�_�_�_ �_o#o
oGo.oko}o do�oO&O�o�o�o 1�oUg�O�� ����L	��-� ?�&�c�J��������� ����ڏ���;��o �o~��������˟ݟ 0��t%�7�I�[�m� �柣�����ٯ���� ���3��W�>�{��� t�����տ�Z�l�� /�A�S�e�w�ʿ��� ����������+ߒ� O�6�s�Zߗߩߐ��� �������'��K�]� D����Ϸ������� ���d�5�G���k�}� ��������,����� C*gy`� ����������}�,ew����)S�W��/ "/4/F/X/j/��/u/ �/�/�/�/�/?�/0? B?)?f?M?�?�?�?�?�Q�����$UI_�POSTYPE � ���� 	 �?#O�2Q�UICKMEN � KO&O�0R�ESTORE 1�6��  O��?X��O�C�OX�m�O�O__ '_9_�O]_o_�_�_�_ H_�_�_�_�_o�Oo 0oBo�_}o�o�o�o�o ho�o�o1C�o gy���Zo�� �R�-�?�Q�c�� ��������Ϗr��� �)�;����Z�l�ޏ ����˟ݟ����%� 7�I�[�m�������� ǯٯ�����
�|�E� W�i�{���0���ÿտ ���Ϯ�/�A�S�eϼw�1GSCREA@?�FMu1s]c�@u2��3��U4��5��6��7��y8���2USER��d�ϫ�T����ks�ê�4�5�6�7��8��0NDO_?CFG 7K<�;�0PDATE �������ޝ4B��_INF/O 18����RA0%}���Q������� �'�
�K�]�@��d� �����������*L���OFFSET ;FM�Ë@ � b�t������������� ��N�UL^� ������&VO�(
L*�UFR�AME  ��d֑�RTOL_A�BRTp�ӈEN�B��GRP 1�<�IRACz  A������	//-/?&I/[/�@@�U�iѠMSK � ��ӢNm�%��%��/�_EVN��$c�
6Uҫ2=I9hi��UEV�!t�d:\event?_user\�/T0#C7Y?)�F�<L1�SPR1W7spo�tweld�=!�C6�?�?�?�@�$! �/h?&O[OGl�OJO 8O�O�OnO�O�O�O_ �O�O�Oe__�_4_F_ |_�_�_�_�_�_�_=o ,oaooo�oBo�o�o xo�o�o'�o�j)6?WRK 2>@�8#8"�� y� ���
��.�@�� d�v�Q�������Џ� �����<�N�)�_�������$VCCMfU�?\ݨ�MR�2E8;<�"��	j���~XC�56 *�����h� �5�i�A�@7 p? ȗ� 	;[�e�Ȇ����ů����^�9%A���ٯ*�� B���E��I� ѯj�����]�����ֿ �������0χ��fπQ�cϜ�O����ϥ�I�SIONTMOU�? ��ů�FU��U�(� FR:\���\u�A�?  �߀ MC*�LO�G7�   UD�1*�EX[�E!'� B@ �� ��o�r���o������d� �  =	 �1- n6 � -����Ҭ6,x�ր�1�=���:����n�P�TRAIN����1�E!�A�d��͓G8; ( ��:��S��������� ��-��1�?�Q�c�u��������T���_��R�E��H�����LE�XE��I8;�1-�e��VMPHASOE  ���A����RTD_FIL�TER 2J8; ��R���� ���1C#� �t��������//��SHIFmT�"1K8=<���/p/3��O/u/�/ �/�/�/�/�/?�/? )?b?9?K?�?o?�?�?��?	LIVE/�SNAP�3vs�fliv4�?�}�� SETU�0BmenuOO�?`}O�OfB/%L���	|H{O�O��?�J�� �@-�AdB8�����K�M�QR�S����	'-G_ME�0�ļ�/!kMOM �zWq�WAITDINE�ND����TOK�  噰\���_S��_�YTIM����
lG�_,m�_Ok�_�/j�_/jo�XRELEK_g���Q��֗Q_ACT�0^h(q�X�_3� N��)r%��O_��rRDIS��0�n�$XVR��BO �$ZAB�C͒1P�� ,����2g7ZIP
�CQ����/�A�S���zMPCF_G 1R�J�0��w��a�MP�sS���<������8����v�4���?�  �������������m��Da��q~D�Q����?��\��*�X>�<����A���#c>�C�~���"�4�;B� T�f�v�e�Ο�����A�2�6���´ $�6�>Ȇ�n�h�z��� ��ȫ�pt��T|��w��YLINDqU�|�  �e� ,(  *)�:���&�0c�J���n� ��� Ͽ�#��s�(��!� ^ϡ��ϔϦ����e� K� ���$��y�Z�l���{��2V�+q đ����������ߠ��٧�D��ז^�A����SPHERE 2W	�̾Ϛ�� �������<�O�*�<� ��`������}����� ���I�[�8��\ CU�������pZZ�f ��f