��   ��A��*SYST�EM*��V8.3�0340 11�/9/2020 A   ���	�BIN_CF�G_T   X� 	$ENTRI�ES  $QW0FP?NG1FU1O2F2OPz �?CNETG  ��DNSS* �8 7 ABLE�D? $IFAC�E_NUM? $�DBG_LEVE�L�OM_NAM�E !� FT�P_CTRL.{ @� LOG_8	��CMO>$D�NLD_FILT�ER�SUBDI�RCAP� H�O��NT. 4� H�9ADDR�TYP� A H� NGGTHOG��z �+LS/ D �$ROBOTI<G BPEER�� �MASK@MRUv~OMGDEVK�%RCM+ ;$�� ���QSIZNTIM�$STATU�S_�?MAIL�SERV�  $P�LANT� <$L�IN�<$CLU���f<$TOcP7$CC5&FR5&�JEC!�EN�B � ALAR�B�TP�w#��V8 S��$VA5R)M�ONt&���t&APPLt&PAp� u%�s'POR ��_T!["ALER�T5&2URL �}�#ATTAC�[0ERR_THRO�#US29�38ƚ CH- �[4MA�X?WS_1��y1MOD�z1IF� $y2 � (y1�PWD  ; LA�u00�NDq1TR=Y�6DELA�3z0|��1ERSIS�!�2�RO�9CLK��8M� ��0XML|+ �#SGFRM�#�TCP�OU�#P�ING_RE�5OAP�!UF�#[A�C�"u%_B_AUZ�@���B�"COU!�U�MMY1�G2?��RDM*� $GDIS�%J@Io�/ 3 $ARP��)_IPFOW�_��F_IN�FAD� �H{O_� INFO���TELs P�~���� WO�R�1$ACCE�� LV��RF�!βICE�0�Q � �$AS  �����Q��
��
�PV�1m@�W�%���QI0A�L�_�Q'0 �X
�
��F����%Bb;e���� #m��!��Qzo���$ETH_FLTR  �Y�.` �P ���B����k�� #m2�k�RSHAR� 1>#i  Pvo,8dXG|?� c������� B��f�)���M���q� ��䏧��ˏ,��P� �%���I���m�Ο�� 򟵟�(��L��p� 3���W���{�ɯ� �կ6���Z��~�A� S���w�ؿ������ � ���V��z�=Ϟ�a� �υϻ��������@�l�gz _L�11�m_x!1.{�0I���z�1���25c5.�Ղ����@ey�2�ߒ��Ц߸�������3�ߒ�o��0�B�T���4p�������������5���_� � �2�D���6`���@���������������6AMY�(M?Y��p���P� Q� 8�<r����@��%7 �P gy�J���� �	//-/��� Cew/b,Q/��/�/�/��/�}iRCo�nnect: i�rc4//alerts�/9?K?]?o? 5�/�?�?�?�?�?�?��0cP9a�� �?0OBOTOfOxO�O�O��O�O�O�O�O_�$�?3_�`("_[_�/_��_�_�_����`a�i�R>j�U�Q�Q�t)�eI DMZc�an�$TCPIP�[b�mi(`=aE�L`��e�Q��`H�!TB�o�rj3_tpdb/� m�vQ!KC�L�o�kv_.��V!CRT�o�oF`�d!CONSGz�j�asmonL�d