��   ?Q�A��*SYST�EM*��V8.3�0340 11�/9/2020 A   ����MN_MCR�_TABLE �  � $MA�CRO_NAME� %$PRO�G@EPT_IN�DEX  $OPEN_IDa�ASSIGN_T�YPD  qk$MON_NO}�PREV_SUB�y a $USER�_WORK���_�L� MS�*RT�N   &S�OP_T  �� $�EMG�O��RESE�T�MOT|�H�OLl��12��STAR PD�I8G9GAGBzGC�TPDS��REL�&U�s �� �EST�x��SFSP�C���C�C�NB��S)*$8�*$3%)4%)5%)6�%)7%)S�PNS�TRz�"D�  ��$$CLr   O����!������ VERSIO�N�(  ����!IRTU�AL�/�!;LDU�IMT  ���� ���4MAX�DRI� ��5
�4.1 �%� � d%�Open han�d 1����% t?�? �"  1�3�0Close�o?�?�?	O�9�7Relax�?�?GOmO�9�6j82oOPO�OtO�3�?�O�O&_�O �6 +O__�_;_�4�F�_�_�_�_�[�3 ��(@�_6o�_Zo	oo �o?o�o�ouo�o�o�o  �o�oVS�; M�q����.� �R�����7���[� m����ߏ�ǏُN� ��r�!�3�m���i�ޟ �����ß8�J���3� ��/���S�e�گ��ׯ ���ѯF���j��+� ������ֿ����ϻ� 0�߿�+�x�cϜ�K� ]��ρ��ϥϷ���>� ��b��#ߘ�G߼��� }߷���(�����^� �[��C�U���y��� ���$�6�!�Z�	�� ��?���c�u�������  ����Vz); u�q���� @R;�7�[ m���/��N/ �r/!/3/�/�/�/�/ �/�/?�/8?�/�/3? �?k?�?S?e?�?�?�? �?�?�?FO�?jOO+O �OOO�O�O�O�O_�O 0_�O�Of__c_�_K_ ]_�_�_�_�_�_,o>o )oboo#o�oGo�oko }o�o�o(�o�o^ �1C}�y� ��$��H�Z�	�C� ��?���c�u�ꏙ��  �Ϗ�V��z�)�;� ����柕����˟ @���;���s���[� m�⯑����ǯ�N� ��r�!�3���W�̿޿ ��ǿ�ÿ8����n� �kϤ�S�e��ω��� �Ͽ�4�F�1�j��+� ��O���s߅߿���� 0�����f���9�K� ���������,��� P�b��K���G���k� }�������(����^ �1C���� ��$�H�	C �{�cu��/ ��	/V//z/)/;/ �/_/�/�/�/�/?�/ @?�/?v?%?s?�?[? m?�?�?O�?�?<ONO 9OrO!O3O�OWO�O{O �O�O_�O8_�O�On_ _�_A_S_�_�_�_�_ �_�_4o�_XojooSo �oOo�oso�o�o�o�o 0�o�of�9K ������,�� P���K�������k� }�򏡏�ŏ׏�^� ���1�C���g�ܟ� ��ן$�ӟH���	�~� -�{���c�u�ꯙ�� ��ϯD�V�A�z�)�;� ��_�Կ����Ͽ�� @���v�%Ϛ�I�[� ���ϑ�ߵ���<����`�r�!�[�
Send Events��S�SENDEV�NT��Q�.��� %	��Data<�߶�DATA�Q��-��%��Sy�sVar;��SY�SVw���O�%�Get�x�GE�T+����%R�equest M�enu���REQOMENU?���� ]ߞ�Y���}�+����� .��d�7 I�m����* �N����� i{��/��/ \/G/�///A/�/e/�/ �/�/�/"?�/F?�/? |?+?�?�?a?�?�?�? O�?�?BO�??OxO'O 9O�O]O�O�O�O__ _>_�O�Ot_#_�_G_ Y_�_�_�_o�_�_:o �_^oooYo�oUo�o yo�o �o$6�o l�?Q�u� ���2��V��� ������q������� �ˏݏ�d�O���7� I���m�⟑���ݟ*� ٟN������3����� i���𯟯�ïկJ� ��G���/�A���e�ڿ �����"��F���� |�+Ϡ�O�aϛ����� ߻���B���f��'��a߮�]��߁ߓ��$�MACRO_MA�XX�������Ж�SOP�ENBL ���2��ݐѐ��_���"�PDIMS�K�2�<�w�S�U���TPDSB�EX  K��U)�2�����-�