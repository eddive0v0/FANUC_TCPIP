��  �A��*SYST�EM*��V8.3�0340 11�/9/2020 Q  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  �  �ALRM_�RECOV� � � ALM"EN5B��&ON&! �MDG/ 0 �$DEBUG1PAI"dR$3AO� �TYPE �9!_�IF� ` �$ENABL@�$L� P d�#Uژ%Kx!MA�$iLI"�
� OG��f �%CAUSOd�!PPINFOE�Q/ �L A� �!�%/ H� �'�)EQU�IP 20N�AMr �72_O�VR�$VER�SI3 ��!COU�PLED� $�!PP_� CES( C p71s!Z3> ��! � $�SOFT�T_I�D{2TOTAL_�EQs $�0�0N�O�2U SPI_I�NDE]�5X{2S�CREEN_84no2SIGU0o?|�;�0PK_FI� �	$THKY�-GPANE�4 ~� DUMMY1d�TDd!_E4\A!R��!R�	 � �$TIT�!$I��N �Dd�Dd �DTs@�D5�F6�F7�F8�F9�G0�G�GZA��E�GrA�E�G1�G1
�G1�G1�G �@!�SBN_CF>"
� 8F CNV_J� ; �"�!_CMN�T�$FLAGyS]�CHEC��8 � ELLSET�UP � $�HOC0IO@� }%�SMACRO�ROREPR�X� D+`�0��R{�UHM�P�MN�B�! UT�OBACKU��0 �)DE7VIC�CTI:0�A� �0�#�/`B�S�$INTERVA�LO#ISP_UN9I�o`_DO^f7��iFR_F�0AI�NA���1+c�C�_WA�d'a�jOF�F__0N�DEL��hL� _aAqQbc?Yap.C?�Y`�A-E��#%sATB��d��AW{pT $DB� g"� =S�$MO�0B x!kq� \� ;VE~a$FN!�p�d�_�t�rdTM�P1_F�u2�w1�_~c�r~b MO<� �cE D [�mp�a���REV��BIL0�!XI�� �R  �� OD�PT�$NOnPM��I�b�/"_�� m�蘁H��0DpS �p E RD_E�L�cq$FSSB�n&$CHKBD_YS�r�aAG G�"$SLOT_�H�2��� Vt�%��x�3 +a_EDIm   � �"���PS�`84%$�EP�1�1$OP��0�2qc�_OK8ʂ� e0P_C� c��+dR�U �PLACI4!�Q���( �a�p9M� <0$D������0pB�UOgB,�IG�ALLOW� �(K�"82�0VAaR��@�2�sBL�0;OU7� ,yq�`�7��PS�`�0M_Ox]d���CF��7 X0GR`0�z�M]qNFLI�<���0UIRE��$ށwITCH�sAX�_N�PSs"CF_�LIM�t=�SPEED�!���P��p�PJdV���u�u�3z`�P6��ELBOF� �W��W�pH� ���3P�� FB ���1��r1���G� �� WARNM�`d܁�P����NST� CORz-PbFLTR۵/TRAT�PT `� $ACCQa�N �r�pI�o"���RT�P_S�r C�HG@I�Z�T(���1�IE�T�Y1�݀�� x pi#�Qʂ�HDRBQJ; #C��2��3��U4��5��6��7��U8��9s!k�M$��	3 @F TR�Q��$�V����C�FN�_U�pY�k�OpT <F �������#�I2q�LLEC7�>"MULTI�b�"��A!cj DET_��R  4F S�TY�"b�=*�)�2��o���pT �|� �&$L�>�+�0�P��u�!TO���E`�EXT�יၑ8B���"2����
�t k0F�RLƯ�r�q���� !D" �M��Qm� �蠋c������"��G�1�ց�qM���P��! �����# L0	����P �pA��$JO�B,�ǰR�0�TRIG��$ d������ �� �K� l��弧Ҹ`�0b% t��F̝ CNG0A�qBA � ��x��
�!v�� � ��z�0�P{`�,R·&ΰf�PtЎa�!��"J!�_R��rCJ$�(J)�D�%CHӽ���z@h�P�Z�@ '�.�RO`�&�סIyT�c�NOM_�`����Sj��pT("�@�݉��P�ǭ��RA�0�2&"��>�
$TFV w�MKD3�T���`UC1�[�g�'�Hgb�s1q*E���\Ѕs�qŦpgAŦsA�YNT�q��P|pDEF�!)��G�PU8/@�܌���AX��Ģ�eT;AI~cBUFņ�||psQ* � �'��PI�)�P�\7M[8Mh9� k6F>\7SIMQS)@wKEE�3PATѠ�"�%"�"$#�"�L6�4FIXsQ+ �L��AdC_v����2�3�CCIh��5PC9H�P�2ADD�6,A@E,AG,A!H�_�0�0_,@�foA)�Ԁ zFK� '�=$#�"��4E��, l���7zp F�CE�C!F+HS@�EDIS�G�3�-�P=��MARG���r�%�FAC
��rSLEW<���x;�M��MCY.����pJB����
aC�Wv�p�U҅�X/ �?��CHNS_EMP���$GE g݀_�} ����pP�|!TC9f��y#a���NdW#�%I��r<��<�JR|�И�SEGFRoP�IOj�ST`�L3IN׃�cPV����!�$0�����b'��b�B��1` +`��	��a	`���a��Pܠ��At��Py�QSCIZ���ltKvTVs0E pz�y�aRS%Ѽ� uc@Q{k�|�`�xZ`�`�Ld�| `�vCRC ɥ��!����t�`%�9a8˭9b��MINQ�9aP7��q�D�YCk�Cz��le��50�p ���EV���Fˁ_
leF��N����Q۶��X%+4,��#=0|!VSCA�} �AY��c1G"�2 �>�
/Ψ`_rU@�+�@w][��i %�7�"�}R��3� �ߠ�߱���5ġR�HwANC��$LG��l�*1$�0ND�סAR�0NK�a�q��acm�ME�1��n��A0h�RA��m�AZ�����X%O`�FCAT���7`�vS�P.
ADI�O��� u��pWP ������ⁱGv�BMP�d�p�D&ah�AES�f@̓�W_P�BA�Sk�s��4  ��I�T�CSXh@�w�5��	$�K1�T��?sCb��Ny`�aBP_HEIsGH71��WID�06�aVT�AC��u��!AQP0� �\�EXqP+�L�@��CU�0_MMENU��6��TIT�1	�%���a�!A1ERRL���7 \���q��sOR�D��_IDG�=�QUN_Od��P$SYS���4��j��Iϡ	�EVG#|�a��BPXWO��z��8��$SK��*2�QDBT(�TR�L��9 �� AC�`�u䈠IND� DIJ�4 _Z�*1KԬ*�W�PL�A�RWA.�tТSD�A�ת!��r@Y�UMMY9�ª�10���¾���:	�A1PR�q; 
��POSr��g; ��[$S$�q�PL��<��H�S@��=�'�C��>4�'�ENE�@T�{�?S�S��RE�COR.�@H ��O�@;$L��<$��62����`�_q�b��_D9�W0R	Ox@�aT[���b��.�F��������PA�c���bETURN,�V�MR��U� ��;CR��EWM�bmA�GNAL� 72$L�A�e��=$P��>$P٠= ?y�A<�C���@�DO�`����:���GO_AW ��M�O�a)�o���CS�S_CNSTCY�@A L� ^�C`'� ID[^�2
2
N��O���ـ}I�� B PNPfRB^rzCPI{POvI_BY�R�}�T�r��HND=G.�C H�DQ�kSP�s*�SBLI�O�F��0��L�S�D��0N0�	FB��FE��Ch��жE�DO&a-sO�MC`{�4(�C�rH��WFPB����SLA�P�F�bIN� �N3������G� $$ ���P]��v��v�ޕ����!o�"��#I!D�&L�&W�";$gNTV*3"VE 4��SKI��as�3�'2�b&aJ�&aM��mdSAFE,d�'_�SV��EXCLUt7ѻ���ONL`��#YcL���4��I�_V8���PPLY�y�R��H[0'3_�M@�NPVRFYI_S�2MS�O@���k6�1�~3�#O�t !5LS�E��35H�£1�`%�P���$��t5�%� Hy��TA2�DP��� �_SG�� I � 
$CURB�_�
�B �������#H��3F��UNM��DZD@���l�{IxA��JZ�F ��EF��IM�J @F]Bk��pOTb�k�ԋѭ5��h�P�и@M� NI��!K��
RwPA!(T�DAY��LOAD�j��R�ӵ2 �E�F/�XILy�Ĉq}�OhPe�D�_RwTRQ�QM DF����P�r�S`�ThU 2L�`���Qkp�P���Q�QN 0�A��QA�t�R���DUtb���"�CAB�a�O�B�NS�QW`ID�`PW���U/q� �VjV_�P�P����DIAG�1�aP�� 1$Vb�HuT�l��u�t� �j���rR�p�DQ�tVE��Y@SW�ad�p7`q�d�U�PM�p�QOH�Uf�QPP�`�sIR���rB��Fb�S��q��q �@3r��-x ��-uj�#e�PO��P���uR7QDWuMS���u�A�u�b�tLIFAEZ��C�p���rN�q �r�uxA�s�rI�xB�Cp���NC�Y���r�FLAW�y@O�V���vHE'ArSOUPPO2���rbS�_E�)E�_Xf�(h���s�Zp�Wp�p�`s���xA���XZ�����qY2ˈC
�T������eN됕exAJJ� v_��q���/���Q `[ CA�CHE��3�SIZ��v*��"j�N� UFFIo� �p����Ե3��6����Mܞ���R 8�@KE�YIMAG*�TM��ᄣ��D��q�>��OCVIE�`�'S ���Ll$@)#?� 	��%����T�P�ST� !��`!��@!�VP!�|�0!�EMAILy��1Q��� _FAU�L��U� �9��C�OUz ��T��|aV�< $��zS��PC`IT�#BUF@F�)!F�Oy�o�D�	B��nC($�������SAV�Ţ�`� ��`���|FP
�z���d� _���"P_�#OT�����P[0���� B��AX��-�I����Wc7�_G�s��YSN_$q'�W�RDuTY��#rMb�T��F+�fP^@D�&�X������g�C_��&�K��8�4B�3��R��2�q��D�SP���PCy�I�M�pÖ��#�Æ`U`M�:���K0d�IPm#0�q	�o�TH��=�c�mPT��p�HSD=Im�ABSCz$��o�V� �Я�&�`��QNV�!GO�&ԑ�$mƸ�F�aаdR�����,�SCxbk(�M�ER4�FBCM�P3�ET�1�Y6��FUX�DU���\���%2CDf���z��u��R_NOAU]T�  Z�P4 ��"U�IUPS�Cʵ@�C�1ϱ���㍰��[H *�L t�3���� �@�0�#�����A��@VQ��1�扑��7��8��9���p���1���1��1��1��1���1��1��1 �2R�2���2��2��U2��2��2��2��U2 �3�3��3��B��3��2����3��U3��3 �4� _�sXT�aQ\ < ���I簉���3�FDRxd]T��V�0���r�.�rREM�`F��r�OVMI�>AGT7ROVGDT�gMXvING�fNuaIND��r
�<�а$DG��:s�p��u�aD�VpR�IV���rGEA-RI�IO�eK7�tN�%(hQ�x0h `�>�sZ_MCMÀ�q�;�UR��^ ,<�1? �� s?� �a?�!	E�0�!�����_P}pP���`R�I�դ$�aUP2_� ` VPģTD����3�#?@�!�'�%��%BACܲa T��Ţڠ�A);@OG�.5%�CT����IF�Iq���x�:pC5PuTV�MR2
�b �3LI��3#/5/�G/^|��u7_�D��R_�A�԰`M�|/-DGCLFuoDGDY_HLD�!��5�v��tz3�c��P�9 T�F9S]��d P� �B��0��а$EX_�A�H�A1kPl���@53[5V�G:�
ge ����SW�}O�vDEBUG4LWR�eGR� �U�ӷBKU��O1a� pPO�P�YoPع�BUoPMS�0OO����QSM�0E������ _E f� �`Ȱ�TE�RM�Ug�U���O�RIe0�Qh�U���GSM_80Ţ�Pi�U�� �TAij�VD�X�UP�k�s -��f$�U>a`g$SEGfjx@�ELTOV�$U�SE��NFI"���bn �q+�d]dh$UFR02���a����	@OT�gU�TA� ��cNST`P�AT��?��bPTH	J ���E�:��АbART+��e|�+�V�ΏaREL<z9�SH�FT�a q.x_SEHI�M^���f $`��xj)A�0OVR���ǲSHI_p&DUz4� %�AYLO��AֱI�ѻ# qk�%�k�ERV���q�yz ��g`<r4_0&����_0RC�!9�ASY1M	�9��aWJ�g���E�#*qV���aU�z�`ֱ.u|���DuP����pYѪvOR`ML�3Z�GR�Q1Tl��oR�V�`�`A" ��B��m �>�b6.71TOC�a�QT!k�OPZ2���}����303OYߠREM�Rm�9�Oѐ$�reT�R�e��h�Fq�/4e$PWR�I�M���rR_C�#tVcIS`sb�UD�#�fsSVW�B��b �n� $H.56�_�ADDR�H�QG r2�'� �
�R��~�.o H� S��Q��4_���_���_���S�E�A�HS��M�N�Ap `T���_����OL����v���ּPACR�O���aS�ND_C�����qٔZ�ROUIP���_X���@��1��25���?�4  ?�<@���?���?���6�2AC�IO��W��D:���J���1Sq3 $� ;�_D� �P�M���PRM_.�~H��HTTP_��HQar (�OBcJE��"�/4$��LE�c��s � ���AB_��T�SS�S� �D�BGLV��KRL~ÙHITCOU�[BG��LOF�R�TEM�ī�xe�a7�f�SSQ ��JQUERY_FLA��G�HW��aQatZ����F�PUR�IO�h����u�у��ѿ� �IOLN�2u��
@C���$SL�2$INoPUT_�1$��bi�P m�D�SL��Qav��gߢԝ�=�s��=�B_�IO�F_�AS�Bw%0$L :0'�:1�q��U`|p§aTժ�_��pHY�� �����UOP�Ex `��>��� ��hᣐP�Ã��^����x�� U}J	y � � ;NE�wJOG�g��7DIS�3J7���+J8��7!PI�a��>�7_LAB�a3�x�����APHI� �Q��9�D�@J7�J�� �@_KEY� �K�L�MONQaz� $�XR����WAT�CH_� �s98��E�LD.5y� n�E{� ��aV�(���C�TR@s����%R� LG�|���~DSLG_SIZM��� &�@%��%FD0I$;�Q2#�P =/" _�+��@���ЩR ��P��S���� �ťV" ZIP�DU�r��N��3R}J���@P�A��]�"d0U�-�L6,7DAUREA��/�h^GH0������BOO2~� C��ӐIT�Ü>@���REC�SCR�N����D��FR'�MARG�2Ҡ����ӐN�"����S3���Wp���A��JGMG'�MNCH����FNtd�J&Kp'PRGn)�UF|(�p|(FWDv|(HL�)STP|*�V|(e0|(�|(RS"�)H�+��C�t�# y���1P#'G9U籐$@"'�r0&���"G`)�WpPO�7�*��#M�07FOCwP(EX.��TUIn%I�  #�2,#C8#Cl p!��p��v3@���p�N�sANA�҉b�p�VAI��CLE�AR�vDCS_H�I\T�Bu��BO�HO&�GSI�G�HS�H(IGN; ��Mm!���T٤�@DE�(4L1L\�C���BU�PR`����pT4B$F1EM�����)�rRQa����pW��\Ρ4�OS1zU2zU�3zQYT�AR`� ����΁�esԲs�$J`�P�r��O�P���a�VST?�RiY���a �$E�fCkW��&f9f8�U��V�� L���_�#�|p��U���וE���֕YU�_ � �� .�6���c� �MC � =���CLDP?�J�TRQLI�[����i�dFLG���`���srAD��w��LD8utuORG��!2 1r��vyxu��t���dд� ���t"5�du� PT�`��bp�t}�vRCLMC�t`}��y��YPMI������ d)�QRQz����DSTBP���P [��h�AX��bi�k���EXCE�Sy�;�M��U��O��d;��V�5�Z�]�_AW�\���������`KB� q\�����$MB���LI�I�REQU7IRE�cMON�
��a�DEBU��;�L:�`MA� ڰ �Л�����q;�ND
>S��'��ړ3DC�2:IN�7GRSM�����@N����F3��PST� �� 4}�LOCf�VRI���UEX\��ANG�RY�;�ODkAQA�K�$t�1RBMF��]���Y��b0�eǥC�SU�P�eYPFXS�I�GG� � � ���b�wÓc:6�d���%c�?��?�.�<��DATACWk�EE��E�����N"R�� t��MD��I��)���@��-���H�p��ᥴX�!�AN�SW!��`Q�1��D���XQMO�� ���[ ÀCU; V㰘 px���LOj���H��5�W�3�E���tU�M�;�RR2B���� (E�NA��q d$CALIIa��GvA��29��RIN� ��<$R���SW0���)�A�BC��D_J2SqEu�Y���_J3��
��1SP���Y�	P���3�"��Y��J�J�Z՞r�O�!QIM��(�CSKAPz��1oC��Jq(�Q�ܺՠպհ�e��_AZ�rV���ELxQU��OCMPs�)����RT��G�c1���5��P1�9�tf�G�ZE�SMG0�}��Օ`ER������PA �S(���DI��)�JG�`SCLܤ���VEL�aIN8�b@��_BL�@Y����Z�J��������ܭ�IN�ACcR���	"x��
f`_u�!�<��YP�9�܂�F���YPDH褀;����iP$V0����'A$d�b���P`��qy�B���H �$BEL���|�_ACCE��� �����IR�C_����ppNT<�Q�S$PS���bL  ��&s�	x1w@
PATH���_��_3..���_@wQ�� ��rb�CC ���_MG !$D1D���`�FWE�~�`��������DE��PPABN6ROTSPEE�{Q8�`��{QDEFb���~. $USE_��JBCP��C�0BCY����q s�YNA�A��}yм�}MOU&�NG�R� O��Q�INC�m����h����i�ENCS���d�Y�&��f�# I�N�RI.%���N�T����NT23_�U��`�A#LOWL��A~0��`�a&D�a0Y�C���`���C�,�(&MOS�@�M�O�ǀ�wPERC�H  ~#OV��  �'�Q�#F�d"&�F�� 
�gm �@w�A. 5LADw��v�)%�d*�_6z&TRK���QAYI�3쁏1.�5�3�n������PMOM  Bh��sp"�W����a�3azR��DU���S_BCKLSH_C.!E��&� ��-�?D�JJ���CLALBP'"�q�0܀N|ECHK�`�US�RTYJ�N����T:S�eq}�_c�$_UM���IC�C����C(7LMT�_Lwp� ṮWE]&P[P !U,�5A�+0gT&8PC�!8H�`|�d��EC�p�bXT��.�CN_��N���V&�SF���)Vg�a�	'|�Q.
e�XCAT�NSH������ eq
A
&F�/F�Z� 3PA�D�_P�E�3_�`���6� �a�3�d��EJG�p���cO O�G�W��TORQU Y/Ւ#�9� ?��"��� r_W�5�4C��<t��;u��;uIC{I
Q{I��F��.qaҐx,pѽ VC��0b�Z���r1�~���s��uJ�RK�|�r�v�DBҲ�M���M�_D9L��:2GRVBt;�0��;����H_L��b i�COSv��v�LN�p������𛉀d���mq׊Ō�q�Z���&�MY������TH��6�THET=0j%NK23��`�l�㣀CBe�CB��C��AS���mt����e�SB��p�'GTS��(C�m��=�cM��ԃ$DU�@C7����� ���9QF�s�$NE��ؠ�I���C)���T�A�X�����h�s�s�LP!Hv�_�9%_�S�ң Ņңԅ_���������V��V����V�ʪV׫V�V�V*�V�V�H��E��²��?aٸ׫H�H��H�H�H�OJ��O��ONɹ�OʪUO׫O�O�O�O�O�F_������Ņ�Ė�SPBAL�ANCEQԃQLE6͐H_X�SP��9�ņ9�ԆPFUL�C=�d�L�d�ԅ&�1=��UTO_�@�e�T1T2����2N �A��?�Ԗ��1f�D�(5���1TP0O����>,pINSEG��!�REV�փ "!DI�Fy5K�1�0��1� OB&�lAE��7�2p?�A$�LCHgWAR��AB�a~�5$MECH���%����FAX�1P�JT��z���З 
p��q��%ROB� �CR.��R[�M�SK_���� P+ ��_WR��r0�?{41	b4 20�1#JD0���IN���MTCOM_C|�p��  � �8�$NORE�$#���t���� �4�0GRr��FL�A�$XYZ_�DA��nC DEB�U�� ��t�� �0�$uCOD[A� ���2���0�$BUFINDXr2�C MOR#�� H-��0���F�B �0�JD$�����QVPTAA�+�2G6� �� $SIMUL��` 13�3OB�JE;ТADJUyS�� AY_I�A:	8D�OUT�`����0�_FI�=@T+p4 ��X�@3p3�A�5Dr�FRI(CXT8ER�O�` E3q[0�O�PWO�p'�,> SYSBUq�( $SOP��A�yU�3�PRUNv��PAC�D����0_� NR�X�ABx��PP� IMAG[Ai-�G�P�IMY�"$IN,��!#RGOVRDM�� �aP   #`W�L_��0an%�B�PRB5PX�}`QMC_ED/ *�� PPNq�M�"OQ@MY19NQ�M!�SL;�'� x �$OVSL��S;DI{DEX�S�&H�SP1�"V3p�%N1 q�0378�"A<�M!_SETp'��� @�0K2��AAR)I�� 
^6_��j7��1v1�5� �P �<T���`ATU}S@$TRCI�8H%�3BTM�7�1	I��$4NQ�3� '�� D-�E��"�2z�Ev��1!0l@�1EXE�0�A�!B*B��4S3�Z0.��0UP���9A$Y�' XN�N�7�q�$�q�9 ��PG��� $SUB�1��1�1~�3JMPWAI,`P	3�ELOP�����$RCVFA�IL_CH��AR -���Q�P�T�U��R_PL�3DB�TB�a�R�BWD�V��UM�`TIGp�( ��4`TNL(`TjRRm���`
p	1	XQ� E�S�T�R�A�DEFSP�� G� L-���P_�P��SUNI#�7�PbmAR1@��3�_L�AP�1* �@w�&�����`�� "<0��)�T"N�U�KETb(p��r`P^R&� h� ?ARSIZE`��h1��naS� OR�3?FORMAT��TTcCO� ja�EM���d�SUX�2b�LIOR&�  �$��P_SWItu��!�fLLB&���� $BA̙`1�ON9AKPAM��0=y��BAJ5����2r68v��_KGNOW8cNrA�U9A"ߐDx� �PDC�ryPAY�[�t���y��wZ�sL�1��U!�PLCL_$� ! �s,qv�t�b"�vF�yCRP1O�z�2�tES���w�R4��w�tBASeE$�J��W�_J�q
K�mA��fBu�8�r�q�MAX4P�`�AL_ � $��Qh 1q�!��C[�D:�sEfr�J3������ T� PDCK�� ��T"CO_J3�������
�hr���� ����C_YQ�  � �� �D_1
�z2�tD���n�^�x��m�|TIA4��u5��6[�MOMS @��ȓ��ȓ��B�@�AD��억��PUB{R͔�������b#��` I$PI�$�QM�=q �wk�B1�yk���������iqRM�q�!Ħ~A�Ħ�A
��9d5S/PEED�G�b� �E�T��T�EP-��C��Q+�Q�ESAM(�E�����Ep{� m�$��  k�~@Ƕ�P_�ֹm��k�v{��ŵ��,H��ǳIN̚�c�� 1���B�W�.�W�wˏGAMM��1���$GET9" �D�;�u
��LIBRtcA�RI��$HIb@!_=!�0k���Eh ��1A����LW��4� +��X��7���wP���CEUv�[ �0 �I_b�xu�� L�������ȓu��پ�� �$Ј W1���I�0R���D\��kAT��LE@f�=q�1M�7�ୄP_MSWFLTM��SCRsH7�����!���~B�cSV&�P� A �����#S_SAqs$��eCNO;�C�1fB<��� ��K�����S�C���hrǥ��m�D� a��� � ���в�����U!C��������s ��cMJ�� � ���YLi�K���^SJ�|v!6O� K���BK�- ��O	W���9���M$P��p����DHc�"��1~B�`M��~T2� � $-΍$$W� �%ANG"�q� ���� !��5P&��o���(�c�#��X`O"����Zz�`�@� �y�OM��+�(�:�pL�^�p���CON@��U B�;�_�B� | ၰ��ș@&��@& �࡚m'X&��.���*J���`X$$Pma��PM0QU�� �� 8#`QCO�U���QTHYPH�O/� HYS�`ES-r� UE� ��S`�O�d�   $1P�@�Ŋ2UN�0b��@O��  � P��p45�E��C�RRO�GRA�1A2DO�445IT�Ё1F0IwNFO�� %0hg;�1A�aOI�2�� (�SLEQ@���1��0k6E1S��ޝD� 4#`EN�AB"20PTIO�N�C�T̢/G�TCG�CFA� @#`JX$P��<2���RdH�0OBG)�2S_E9D�@  � �{�K�q�3��E)�N9U�G�HAUT�ECOPY�qI0�L���M��N�@�K��PWRUT �BNV@;OU�b$G92DT}aRGADJ��ͽbbX_ �R$P`pV�pVWnXPnX�[�pV�`Pz�N��_�CYC"ZSNSrE�$ ��LGO����NYQ_FREQ0�Wb��a�d23L�p�b�PnQÓb��5�CRE���#��IFl��s3NA��%?d�_G��STATUx' ��*7MAIL���YsIN��$LASTx�a���TELEMA� �GFEASIA����H �b@�1���f;B����I�0����R=q�!� R�rAIB+A��Ex0�V�a 7vW�Cy��1�U8�I0�pd�lvRMS_TRs��@��sr�7�z��aktB�R��/ 	�b 2� =�_+��ve��w �r� �fe��c�G�'DOUa3;�NHC�R�PR	 @��2GR�ID�1+CBARS���TYC�ROTO\㐾�� %1_[d�!�P��B�OxD�� � �0�PO�Ra3��[���SRV�_`)˄ÆDI�T�^���������4���5��6��7��8���QF��A�#0$VALURs���d��q_�D�� E��u1��aa��=@#AN�㉒qaR�@a>��TOTAL��1���PW�SIJ���R�EGEN����#X�xxI3e%!��� TR^s0���_S��^����CVnQ�D��B8rE��cN��!��42�@ÓV_Hk�DA�~���GS_Y
�rfS��{AR�2� <RIG_SE�ch�Â2�e_80��C_v�`��ENHANC�!'� p�qEqb�Î��INT��� F<.3MASK��ipOVR�#P� N��@`a
�_�*6^�M��Bp[��f8��SLG��>��� \ ��e�H ���Sq�dDE�U��*7Ő�%�2�U�Q�TEj  � (7��҆��J϶�"cIL_M`!d��P㈠�TQ� ��Ë1rpj�eV��CF��P_��op��M��[V1��V1��2�U2��3�3��4�4���ᄠ��������s��IN��VIB�� �İ����2��2���3��3��4��4 �ؾ���#"�������`%��׌ՠՌ�PLv`gTOR� ��INb�p�����  �p���MC_F� 	�B��L����B�ڐM�1IB���#� 1 ��)���KEEP__HNADD��!��$<p��C�_`�䂁��H ��O�!��P��p����G���REM���쑥�;�R�W�U�[de��HPWD w ��SBMo�*��G�1�2�� ~H COLLABu���a������ؑEb�0IT���0��7� ,� FLbq�$SYN��M�C��d�UP_�DLY��#2DE�LAJ �nbY� A�D��PQSK;IP�� Ļ�60aODD���t P_60 _2�g0^ ����	 	Q�	��	%��
2��
@?��
L��
Y��
9�QO�J2R�P��CEX]pT�SY��X�]P��Y�1���PRD�C��b�� ��@ReCg�R4ae��"d�ԇRGEr@sl�:�FcLG�!Pa�SW�IΨ�SPC�3�QUM�_Yt�2TH2N�&�# L 1�� �EF�@11�!� l�����C��AT4�ET1��7 s"k0o4j!�@Y�j!<3\�HOME�"�P<$2D"�J/\/n/�/�/�/�'3D"��/�/�/P�/?!?�'4D"�D?@V?h?z?�?�?�'5D"��?�?�?�?	OO�'6D"�>OPObOtO�O�O�'7D"ֻO�O�OP�O__�'8D"�8_@J_\_n_�_�_�%S��
�1�9 �q=#$��i�S�E��ٷ�a�LbݖJcIOq��jiI�P��GbPO{WE��� 4`� wGbה ۼ�b$DSB�G#NABqՔE C) ����S232Peܓ ���U�P�I'CEUQrt�E3 ���PARITáՑO�PB��FLOW�TR`�c�3����CU+pM��UXT�n���U�ERFAC�tC�Uѐ�cC�H�q� t����_�p��$����O)M۠9�A�T>���UPD�A#�`T�+`҃*�� �x�s!ƞ�FA������RS�PqpQ��� !>�X$USA ��l�Y�EXmpIO6�$�pU�YE��b_�ª�B�#q`�WRp��_�Y�D�����VFRI�END���UFR�AMδ��TOOL�ȆMYH����LE�NGTH_VTE⮄I���[�$S�E�`��UFINV�_�@�5aRGI:���ITI����XX�	�J�G2J�G�1T�U�D�d�u���_Â#O_p�py�၈���n�C	�zŔ�Cp ���ʖ �G��|zr2�� @ 9� qC���d�wu��ysF�� ���p��X� #�E_M�pCT^�H��f��<u6�J	�G#WV�z�G�z��Dh LOCK~��U� ������$� 2���~�D R��1���2��2�3��3���:����@V��V=�"�=�F�V�Ӂ!Ѕ�/������p��xṿ����Pr@ƻ���������E��`����!��AC�CPRs�!�}�S����`�����a�# 0 5�ؠ�V���ؠ���	������
zM�S��� ح��R�qda��$RU�NN�`AX2q��A⸀L�+"��THI�Cx� w �u��F�ERENg���IF��x���I����V��G1&�*Ԅ�1ٲ[��I�_JFR�PR���
��RV_DA;TA�q� RD�Z[ 
�AL� �xՑ �b{�  2� �S�~�`�	� �$ zZ"GROU���!TOT����DS}P��JOGLIYsN�E_P�PrO���\7`��bvK�p_M#IR�.䎐MQ�O�APp��E<�o��t���SYSE�ib��PG��BRK���v$ wAXIa  �������Ҽ�A����H�OBSOC��T�N�����16�$SV�1�DE_OPNsS�FSPD_OVR�4 ����D� �OIR+��PN�P,�F��l,��OV�SFa���d�$�F}�ja2㒓8��ҁibLCHH\RECOV�n���WE�M����RO�Ns���_���� 9@�9�VER��n��OFS9�C�Я�WDE���A����Rh���TRBq6aY�E_�FDOh�MB_CiMkS B��BL��.�u��8�V摁��p���]�Gv��AM���i ������_M�� [r�ec T$C�A��D��HcBK�q�vIO��q,�a��PPA �L1\D��bDVC_DB<���q �b���ja�1���3���ATIO"i`jqcp�U�� �efCAB�����J� �������__p�v?SUBCPU�b�Sv��`_��p"�`'�}���b"�$HW�_C� Ip���'ɣA�x����$UNIT��� � ATTR�I���"�CYCL���NECA�Y�F�LTR_2_FI`#��h��f��LP$���_SCT��F�_�'F_�,E2�*FqS�a��"CHA���-7�1�Pr�2RSD�  �b�����a�`_T��PRO�MFpE%M	`_���Ts2��� s2���5DI�&��tRAILAC4���M��LO�����5��������+PR�S̑{�dA�C�p	��FUN9C!��RIN됫�0|�@�DEqRA�@��� �C7`�CW3ARB�	BLƑ�G��DA�K�!�H�HDA`��AX�C�ELD�p �@S���A�@S�TI��`U�ѓ�$�<�RIA�q�bAF
Q P=��S��U �8���3MOI� P�DF_ꀔ��qHpL�M�FAE�HRD]Y]�ORGEPH�0���|� P�UMULS�E���`'���0J�(�JC�X�S�FAN?_ALMLVBs_a�WRNfeHARD����v�䐟p�@2$?SHADOW��0Ѐ�a�b��_`+q�ї�_,���vAU�Rx4\r?TO_SBR��e����j� ��A	sMPINF���!t6Q�'sREG���aDG�BP��V�p.�l�FL4�%!���DAՀ_X�P�CM��NЍY�B�V  ��� ]���$N��$Z�� �Ҭ����o� �|�EGK�����qAR��#���2?��wP��AXE���ROB��RED���WD���_F���S�Y��!���h�Sr�W�RIE��v� STRP���`��7�E�!�����a��B�����@CD� OTO7q����ARY����.A����#�FI��9�$LINK�Q����y�_���6���8�XYZ�bB�7NP�OFF
 �7�J+��B��yB��0���0}@��FI� ��Є���yB
�_J ��5�����`Ȅҋ8��H�TB�b��C0x�DU �9.AETURa`XgSW����rX���FL�z���#�pu�Y���3x\��� 1��%K�M����31�DBp`%��`'2ORQ�6 �ѳC��}�DB��>��P���%�����\q:�OV	EA���M90=ѻs[� �s[��rZ��`X��aY� � X�O�~@91�P��B� F����=�S�B�_��0�s����ER�A�	EBE��� QC"�Aб�����E�2��Q&QAX���Q�  �!�|�A��+a��� ��@@��O���n������N���1����`�� `��`��`��`�� `��`��`��`��!��� �Rg�DEBU�#$�A�c�2��3�ABGE�;�9V�" 
�Ҷ ���z!$�
�$��$� @A$�O�$�n�$��$��N��T#��R����LA�B���� �GR�O0��l� B_ �1	ƞ�>��`���p����a	�ANDà�E ��<���aF�  ��q��Z�Qi�� ;�#NTq`�cR�C�1=��
��� �pE�RVE���p� $�q��@A�a!��PO�`X �����Q��p�  $.��TRQm�
��Q�2����R2�oP~@_ � l=����fERRҒ�I�V����gTOQ����L%��Ď�z�0G��%%�"��?�!P � ,��2 �뺱RA� 2'� d�D� 7 �p$O��2��PvµOCQ� ��  YCOU�NT���FZN_wCFG��� 4� ^v2T�d�"���m �W k!E�s� ��M�08b�����X��0�FA~P���V�XA������0����O A�P�b�pH�ELkpN�� 5ސB_BASN�#RSR]vm@;��S�!YQB 1�B 2�e*3e*4e*5e*6�e*7e*8�5!ROaOGP� �:�NL�q�)�AB��@C AC-K�INT80�s�U�``x1�)_PUXA��b�2OU��P�@�^x"#�y0��b�TPFWD_KARlLfpZRE���PP��&Q�@QUE]zRO B�2����`�aIb`��"#8�$C0Bv8�SE�Mա�6�`A�S�TY4SO�0�dD�I1�@r�1aǿQ_�TM�sMANRQ�AF8�END�d$�KEYSWITCaHS3h1#A�4HE2��BEATM�cPE��pLEks1���HU�g3F�4h2S(DDO/_HOM�PO�a� EF"�PR���rS�����v�@OaX �O�V_M���`pPIOcCM$��7��v##HK�q� D5�$_w�U�b�2M�p�4�4�%�FORCcsWkAR�R9WOM�p � @��˓�`UU��P�1�V2�V�3�V4�)�O�x0L�R��^xUN�LO.0�ddED��a  �$$C�LASS `����.a�p�7`#`Sܘ0+h���?aIRT?�,o>`�AAVM��K 2� je �0  �5�5a�o�h�o�m �l	�m�pk`!��o2v7u�lV}�b�ah���t{`B�S4�� 1Li�? <�� � �2�D�V�h�z��� ����ԏ���
�� .�@�R�d�v������� ��П�����*�<� N�`�r���������̯ ޯ���&�8�J�\� n���������ȿڿ�h����rC`�AX��� `Ė�s9�%�INf.��<�$�PR�0�XEQ�}�`�_UIPMIl�ja{`L�P�R ji`��tL�MDG �g��`��PIF �k`d��0�B�T߀b�߅ߗߩ߻���, 
���n��o� 0�B�T�g�x��������yNGTOL � �{�pA   ���
�{`Pd�O �� ��=�O�a�s�6b� ��u���2b ������������& J4Z������ ����*<�N`r��zPPLwICA�1 ?je�}����H�andlingT�ool � 
�V8.30P/5�8��
883340��F0!��755�����7DC3������ޝ�FR�A� 6*- s !�� TIVqŔ�>��#UPn1 ���\�PAPGAP�ONf`�.za� OUPLED 1�i� /03?E?W?��_CUREQ 1M�k  P�a7a<��n�?�d}��33b{9b ��Ƨ4H�522�:HTTHKY�?Kx�? �?ZO�?6OHOfOlO~O �O�O�O�O�O�O�OV_  _2_D_b_h_z_�_�_ �_�_�_�_�_Roo.o @o^odovo�o�o�o�o �o�o�oN*<Z `r������ �J��&�8�V�\�n� ��������ȏڏ�F� �"�4�R�X�j�|��� ����ğ֟�B��� 0�N�T�f�x������� ��ү�>���,�J� P�b�t���������ο �:���(�F�L�^� pςϔϦϸ�����6�  ��$�B�H�Z�l�~�0�ߢ��6s5TO��/��#DO_CLEA�N�/q46�NM  �� a?��������g>DSPDgRYR=�p5HI� `�@q�8�J�\�n��� ��������������m8MAX�����17.X�-!*2-!�"PLUGG0�*3��%PRC��B^�"b�'��O���^q4SEGF� K� ��^�p�8J\n8���LAP�( �3���
//./@/�R/d/v/�/�/�/�#T�OTALPy	�#U�SENU"; ��8?�2s0RGDI_SPMMC� o1�C�@@@q2"4O��5 3_STRING 1	�+�
�M� S��*
�1_ITE;M1�6  n�-�? �?�?�?�?OO'O9O KO]OoO�O�O�O�O�O��O�O�OI/O SIGNAL�5�Tryout� Mode�5I�np?PSimul�ated�1Ou�tQ\OVER�R� = 100��2In cyc�lEU�1Prog� Abor[S�1~;TStatus�3�	Heartbe�at�7MH F�aul�W�SAler�Y_ oo$o6oHo�Zolo~o�o�o  �;�?�o�o );M_q��� ������%�7��oWOR� �;o��o I�������͏ߏ�� �'�9�K�]�o�����य़��ɟ۟�PO �;�Q�����6�H�Z� l�~�������Ưد� ��� �2�D�V�h�z����DEV���*� ��޿���&�8�J� \�nπϒϤ϶�����������"�4�PALT�m[ч�5߃ߕ� �߹���������%� 7�I�[�m�������I�GRI3 �;�� s���'�9�K�]�o��� ���������������#5GYk��� R �m��}��� %7I[m� ������/�PREG_�H �!/ o/�/�/�/�/�/�/�/ �/?#?5?G?Y?k?}?��?�?�?]�$AR�G_o�D ?	�����1��  	$�V	[
H]
G��W+I�0SBN_C�ONFIG 
��;IQHRCACI�I_SAVE  �ThA_B�0TC�ELLSETUP� �:%  O�ME_IO]\%?MOV_H�@�O��OREP�_�:U�TOBACK�A�SMFRA:\5+ _5&�@�'`�P5'dReC{� q^ ,H 5-�_�_�_�_�_*o]T���0oXojo|o�o �o�o5%Eo�o�o &8�o\n��� ��S���"�4� F��j�|�������ď�֏��  PQSY�SUIF.SV ���R TL.TM�P DATE.D�^��0�B�T�f�-SI�NI^�5$[E~-SMESSAGw@����A�0��ODE_!D�@zFDV��O��ǟ�-SPAUS'� !���; ((O �2�1��Q�?�u�c� ���������������;�I����TSK�  
�d_j�0PUgPDT����d���ԖXWZD_ENqB��WJ��STA����1���1WSM_C5FO@�5]E�7~�GRP 2�� 	BB�  A܊��9XISI@UN�T 2j��C � 	z���A���Ϭ� ����	���-��=�c�nf�MET� 2u��PNߧ�J���^�SC[RD�1��P	�EB��$�6�H� Z�l�~�]_5*Q{I� ��������(���L� ��p�����������1�k��73QGRn���蟾	UP_NA�@��;	3T_ED���1�
 �%�-BCKEDT�-���J��U /DdD�@-3Sz5*,B�&o�Fs&  ��2�K�wʹ �E��	�-3�X5/|�/|/ ��k/�4�/$/ ?H/��/H?�/�/7?�/5�?�/�??���?O[?m?O�?6 LO�?�O�?�uO�O'O9O�O]O7_�Oe_ �O�A_�_�O_�_)_B8�_�1o���oxo�_�_go�_9�o o�oDo��oD`�o�o3�oCR S_���]��Ug���	 V NO_D�EL'GE_U�NUSE%IG�ALLOW 1z9	��(*��TEM*��	$SERV*¯�Ȁ�7REGх$�܎ȀNUM���	��PMUt���L�AY�Я�P�MPAL��J�CY'C10U�h�R�V���ULSUH�
�j���ӃL��ݔBO�XORI��CUR�_ʐ	�PMCNmVD�ʐ10~�>0�T4DLIȰß<�ˋ$MRߎ�&�&�ϲ����̯ޯ����y	 LAL_?OUT k���(WD_ABOR�o���m�ITR_�RTN�����m�N�ONSTOM ��� ԸCE_RIAS_I������˰�F��U�c����_LIM߂2�` �  N���Nϯ�<��m�`����� ?Ϡϲ���¯�
����p��PA�RAMGP 1U��Ύ�O�a�|s�2�C>  CV����f��z�ߵߗЇ��Б�Ж�Р�Ъ�д�Ԛ٢����������C���ǀ C�ї��+���?��ɲHEC�ONFI��w�E�G_P�1U� 49�� ������������E��KPAUS�19� ,�uG�Y� C�}�g����������� ����1U?e�!�M��NFO �1(�� �=���� �	�����@������%^���ϺA�f��� �D��D�q}�D�Q�6��p���� ˰O����ǩ�COLL�ECT_�(��pEN`���\�nINDEx(����!�1234?567890�� ������H,��)'/L/�|&/8/�/�{ j/|/�/�/�/�/?�/ �/?e?0?B?T?�?x? �?�?�?�?�?�?=OO O,O�OPObOtO�O�Ot�"� � �>�IO "�����O_a_s_�_W[TR�2#](�b8Y
�O�^P�$,]x�Z��Y_MOR"�%� �9�Fe�Fi ^oLo�opo�o�kb�"#�&-mB�?>�>�H���a�Kt�A��PM(���a�-=�Oas�ϗ������^@
����` *cؗPDBO*���Ecpmidbg�C���U�:��qi)��p/���S�  ��e�-�̏�����x��v������7��g�^�)� E��fM���w��>�@ud1:˟����Z�DEF )�o7S)ߑc�b?uf.txt��M�� �p_L64FIX +�Q��� ˓�د��ɯ��2� D�#�h�z�Y������� Կ�ſ
��.�f�x�__E ,� ̀l�~ϐϢϴ���p�I�M�C-�]��6���>���=L�͖��MC&c.�Sd(F�'�%d/5ݤ`t��v��B!!������@�߹���>�T��g1�\�D�y**�~***�}��`U�kx*��CÇЩ���BDw�4��	��a�Ee�3Ec���Et� F��3E�ŚF��B��F���F��YfF�% G��� G	ڳH��3�y?�  �>�33 ;����a�v  nf��q@��a5����b�pA8�a�t�<#�eDQ���7���F�RSMO?FST '�f�VG�T1#`DZ�2!��
�*;��0�R�L�?����<�M��TES�T�0��FRz3hSMx�C�A�z��*e���| C6��B��C�ns���*:d�b�2Iy4<2T�_�PROG �,k%^�/%PNU?SER  �1���KEY_TBOL  -e1]��(��	
�� �!"#$%&'()*+,-./��:;<=>?@A�BC�GHIJK�LMNOPQRS�TUVWXYZ[�\]^_`abc�defghijk�lmnopqrs�tuvwxyz{�|}~������������������������������������������������������������������������������͓���������������������������������耇����������������������A� LCK#D�#STATi/0_AUTO_DOG�����+INDT_ENB�/ �"��/�&T2�/6STO�P�/�"SXC� �25K�p8
S�ONY XC-5�6Q{��p�@���͞b �P���X5HR50��z-tx?�><��?�A�ff�:�O"O  �?GOYO4O}O�OjO�O �O�O�O�O�O_1__�U_g_�\TRL� L�ET��	4 �)T�_SCREEN �-jkcs���PU0MMEN�U 16� <O\�o�u�_oIo ��&oLo�o\ono�o�o �o�o�o�o 9" oFX�|��� ��#���Y�0�B� h���x���׏����� ����U�,�>���b� t�������П	���� ?��(�u�L�^����� �����ʯܯ)� �� 8�q�H�Z���~���ݿ ��ƿ�%����[�2� Dϑ�h�zϠ��ϰ�����b��S_MANU�AL"?�QDBCO�� RIG�Ws)DB�G_ERRL� 	7�[�����ߴ���� O�NUMLIT I���dD
O��PXWORK 18���&�8�J�\�|n�DBTB_�Q� 9<�����K,�DB_AW�AYW���GCP� D=����_AL �/��S�Y!0�UD �H�_q� 1:����0,R0�T�PA�~�6��_M� IS� ���@� ��ONTIM6�W�D�����
2#�MOTNE�ND'"�RECO�RD 1@� y�����G�O�N <����z���G ��Nr'9K ������� ���#/�G/�k/ }/�/�//�/4/�/X/ ??1?C?�/g?�/�? �/�?�?�?�?T?	Ox? O�?QOcOuO�O�?�O O�O>O�O__)_�O�M_8_F_�_�N�ex �_�_�_<_�_�_�_'o�N�U(o_oqo�_��o�o�o�o�NH�I �o�o9$2o�N���p��(������N��_��K�]����TOL�ERENC��B�����L��O�CS�S_CNSTCYw 2A~� h���Џޏ����&� 8�J�`�n����������ȟڟ����"���D�EVICE 2B~� ��r����� ����ϯ����)������HNDGD ;C~�Cz<����LS 2D\� ;�����Ͽ�����=���PARAM CE/���?�)����SLAVE F�~�J�_CFG �G/�)�dMC�:\��L%04dO.CSV(��c��l��A ��CH���n�n�)��=�[��)�-�Z�j�X�W���JPъ�C�_C�RC_OUT �H��<�+ϑ�SG�N I�����\�17-M�AR-25 14�:24��)0=5��6:01���� Ze�7-��)�)�*���o��I�m��P�uG��=��VERSIO�N ��V�3.5.20��E�FLOGIC 1�J% 	���* ������PROG_ENB��.��ULS�� ,P����_ACCLIM^����Ö7�?WRSTJN����)��MO�
���x�INIT K�%
��) v�OP�Tp� ?	����
� 	R575�)���74��6��7R��5��12�����6����TO  ���@���V��DKEXd�d��x��?PATH ���҇A\���I�AG_GRP 2�PI�|O�	 �E7� E?h� D�� C�� C ��B�́�C��nk������C��C�m�B�N�B�zoOB�)�B�k�f3�83 6789012345���B��  A���A���A��A�O�A���A{+As��Aj�RAbJAY% x��@���p��G!��Ae�����B4�h���x�
"�����"�Q�A����A���A����A�� ��hA�x~�Ao�7A�f9X��?$>��mF/X/��h����(�"_�AY�;�AS�TAM�^�AGdZA@��A:bA3%A+�-A$����)�/�/��?�*@��;d�6���@{��@u�-@o��@i�7@c�C�@\�j@Vs{N?\0�5?b?�t?�??@_��@�Z^5@T��@�O�@IG�@�C33@<��@�6�+@/<@(�`J?\?�?�?O�8s�� nE�@h��@b�!@\�0V�ff@Pt@Ihs�@B��@;� bOtO�O�O�O�'6]^_ p_N_�_�_0_z_�_�_ �_�_$o�_�_
olo~o \o�o�o>o�o��C"��!30�2KA�@^>8�Q�r��R?��  *u^7�Ŭ�Fr'Ŭ5AF<Ru^@�p�nv�@�@�pppE�@[ A�h���uC=+�<��
=T���=�O�=���=�<���<��p�q�xG� ��?� �C�  �<(�US� 4rjr�D@����"�A@w�?f�oX� �mf����������ԏ�n��
��.�@��i?�#�
b��\>x�pn�^��G���G�^x���R�����^8�ۑ�5甮��CnB�L�]_u��&�P;�'f�d��aQ{����dD�  D� � C΍��̯ޯ 8����V�ǯPD�ïh������ 3+��Q�ҿ������ ,��P�;�%ZN�Dϥ��CT_CONF_IG Q-��#�c�p�� �STBF_TTSd�
����C�V����MAU^���ҿMSW_CF��R�-  ]z��OCV7IEW�SY�i�����߽������� �G��.�@�R�d�v� ������������ ��*�<�N�`�r����� %����������� 8J\n��!� ����"�F Xj|��/��`��//j�RCR�	T�e&�!�,.V/�/�z/�/�/�/�/�/�S�BL_FAULT� UI*n�1GP�MSK��$7��TD?IAG V��e��2�UD1:� 6789012G345�2��?�P�� �?�?�?�?OO)O;O MO_OqO�O�O�O�O�O��O(� �>�;�
��?%_��TRECPZ?l:
z4l_?��?�_ �_�_�_�_�_oo0o BoTofoxo�o�o�o�o��o�O_/_UMP_OPTION���>*qTRR���!9�KuPME��>Y_�TEMP  ß��3B�Пp�9A�p�tUNI7�����qF�YN_BRK� WY�)8EMG?DI_STA�u&�؟q ��pNC�s1XY� ��o7�*�~y���d ������Ǐ ُ����!�3�E�W� i�{�������ß՟� ���r�,�>�P�b��� �f�������¯ԯ� ��
��.�@�R�d�v� ��������п����� �%�7�I�[�u�ϑ� �ϵ����������!� 3�E�W�i�{ߍߟ߱� ����������/�A� S�m�w������� ������+�=�O�a� s��������������� ���'9Ke�[� ������� #5GYk}�� ����/1/ C/�oy/�/�/�/�/ �/�/�/	??-???Q? c?u?�?�?�?�?�?�? �/O)O;OMOg/qO �O�O�O�O�O�O�O_ _%_7_I_[_m__�_ �_�_�_�_�_Oo!o 3oEo_Oio{o�o�o�o �o�o�o�o/A Sew����� ��_��+�=�WoI� s���������͏ߏ� ��'�9�K�]�o��� ������ɟ۟��� #�5�O�a�k�}����� ��ůׯ�����1� C�U�g�y��������� ӿ���	��-�?�Y� c�uχϙϫϽ����� ����)�;�M�_�q� �ߕߧ߹���E���� �%�7�Q�[�m��� ������������!� 3�E�W�i�{������� ��������/I� Sew����� ��+=Oa s�������� //'/A7/]/o/�/ �/�/�/�/�/�/�/? #?5?G?Y?k?}?�?�? �?�?���?OO�? K/UOgOyO�O�O�O�O �O�O�O	__-_?_Q_ c_u_�_�_�_�_�?�? �_oo)oCOMo_oqo �o�o�o�o�o�o�o %7I[m� ����_���!� ;oE�W�i�{������� ÏՏ�����/�A� S�e�w���������� �����3�%�O�a� s���������ͯ߯� ��'�9�K�]�o��� ������џÿ���� +�=�G�Y�k�}Ϗϡ� ������������1� C�U�g�yߋߝ߯�ɿ ۿ����	��5�?�Q� c�u��������� ����)�;�M�_�q� ������!������� -�7I[m� ������! 3EWi{��� �����/%//A/ S/e/w/�/�/�/�/�/ �/�/??+?=?O?a? s?�?�?�?��?�?�? O/O9OKO]OoO�O �O�O�O�O�O�O�O_ #_5_G_Y_k_}_�_�_ �?�?�_�_�_�_'O1o CoUogoyo�o�o�o�o �o�o�o	-?Q cu���_�_�� ��o)�;�M�_�q� ��������ˏݏ�� �%�7�I�[�m���� ���ǟٟ����!� 3�E�W�i�{������� ïկ�����/�A� S�e�w���������ѿ �����+�=�O�a� sυϗϩϻ������� ��'�9�K�]�o߁� �߭����������� #�5�G�Y�k�}��� ������������1� C�U�g�y����߷��� �������-?Q cu������ �);M_q ���������	 /%/7/I/[/m//�/ �/�/�/�/�/�/?!? 3?E?W?i?{?�?��? �?�?�?/OO/OAO SOeOwO�O�O�O�O�O �O�O__+_=_O_a_ s_�_�?�_�_�_�_�? �_o'o9oKo]ooo�o �o�o�o�o�o�o�o�#5GYk}�_ ��$ENETMO�DE 1Y�U�  �P��P�U��{�pR�ROR_PROG %�z%�V�&���uTABLE  �{oe�w�������rSEV_NUM� �r  ���q���q_AUT�O_ENB  ��u�s�t_NO΁ �Z�{�q�� W *������	��Ā+�*�<�N��HIS���Q�p�_ALM 1[�{� ��T��P+O�˟ݟ���%�rS�_����  �{���rj��pTCP_VER !�z�!�5�$EXTL�OG_REQk�9�ቼ�SIZů���STK����~��TOL  �Q{Dzs��A ��_BWDJ��؆K��ԧ_DI9� \�U��t�Q�rU�STEPa�s��p���OP_DO��qF�ACTORY_T�UNk�d̹DR_?GRP 1]�yށ�d 	e�#��p��x����� �n��So �k� ���W��i�z�d� �ψ��Ϭ�����	�����?�*�c�N�@�� @畱?��߯@Q�j�
 E���R��j��x�d����E7� E??p D����L��D�%��  Cμ��K�B�  ;��  A@E�o�@U�UUc�UUo�&�>�]�>П������E�F@ F�5U��{�L����M��Jk��K�v�H�,_�Hk�{�?�м�Q�9tQv+�8���6h�%7��{�W> O����sO��Gj� ,k��rP�,�FEATURE� ^�UK��q�HandlingTool ��� roduC�hinese D�ictionar�y��LOAD�4D St��ar�d��  NDIF�Analog� I/O��  d� - ��gle �Shift��F �OR��uto S�oftware �Update  � J70 mat�ic Backu�p��art Hg�round Ed�it���708\���amera��F���D pr��nr�RndImM��P�CVL��ommo�n calib �UI q.pc�nf� Moni�tor��wset��tr��Reli�ab	 ��jp �Data Acq�uis����� D?iagnosD������� Docum�ent Viewye���
PC �ual Chec�k Safety�� act.�Enhanced7 UsGFrw ���\weqpxt.� DIO � fi�+ t\j7�e�ndxErr� L�*  � �{s I ��r�� :���T "� FCT�N Menu`v����t I�TPw In�fac%_  48\� G_ �p Mask EKxctg�� o���T Proxy [SvH  5p��igh-Spex�Ski� " #�1��#�mmun�icC ons�apd�!ur ������"conne�ct 2Pdin�� ncr str�u�� I KA�REL Cmd.� LE uaG"t\�ia�%Run-T�i�Env��"K^�el +G sE �S/W�L�icen��[GE�R  �Book�(System)�� R5� MAC�ROs,x"/Of�f� �Pa� MHx�- �: \ac�1�MR� �)��Me�chStopV!t$�  ��0i���Mixx��E ���
� �0od
 wiwtch��Loa� ��4.�6 k G<�1�3OptmUHM �GGW filG� �HF��g�' pmf�O Multi-T�= i�4pa�PCM fun�'{3M"�Po[�D QV^�HRegit0r� �  mpo� Pr�i@F�K _fc�s W g Num Sel�5��� DS� Adju� ����`W
 4 S|XtatuQ/bUC�� �RDM Ro�bot��scov�e�� cctO Rem�0�n���S�ServH10@#CT�XPSNPX� b<2�� "K9<$`Libr���'564@e�� �4H`�ZUSoY0t ss#ag�E�~� "�1n�VVLO�b/I-� pc
�`MIwLIB�mch1o Firm+�8� �b"Acc` hXcTPTX�;��� s Teln�0�m}B����5��4Torqu>
 imula�}n�Tou7@Pa51���m�T_ �QC&�V ev. ocl�eUSB pYoU � iP�a@~WdUSR EVxP�+Unexceptx�P�D{D{f}VC�r�"�"�2�s�VD��j�cV�Hk �uifoV�SP �CSUI�k��XC��6X`Web #Pl�V��9pjăa�+64.f��^ r�>�T�v�
J57�À�vGrid�Qp�lay 76 (���`L&iR;�.t��K�\0ARC; �4 120i��L#AsciiV!eRDAG�d��UplE@��� ޛ@CollW�GuN�� of^QޝPI C  1�s� ��t�0�t8FK���Cy�p � 2*Porie  �ld�aFRL�1a}m͉ RINT��MI DevO0 (&ax2 ,�0�%(}�t\rb�A/��P�asswo��:O�" 64MB DwRAM�

! 0.ڢFRO�qG`��;rciPvis�y6{BW�Welds /cial�4 )���ell���!P�syhK���wmrwd��cXE|�( p�v� w-md�ty	 sPRa���P0�t!1m@.)�8�D�P�����P+�D� 2b a���r�d�r�Pb� q�DrT�1� eged� OL��Sup�r�AR�8sOPT "W� �! � d��; cr�o�V  �SHe[� � ��
gq�<�ues�t;`LO SS��en�tex E��$`p$![b�UsCP�P@ �4YPVir�tW�St�e~�Pd�pn�x��  �� SWIMEoST f� F0��>�ui.�&���ߖ� аߕ�5�1 J����(Fr��ߕ�II)�ߓ�on��!���M!=��	Q�Y���f>�t���mf V��լ���Ҍr��� ?���&P�3��p�Ҭb9���eie����n\p���\R���҂�`A��2�p����!'
!����O����7 J5����5p�ӝ1Q��\ar7����XPR���k "���}��b����`P���lnko����`1��RMJ����;����M�����H54����j883]D#ER�N��Ffh�FM/el���չ1d/ ������d0�/��|B �/�( �/��<��/��9p����.fd�/���ASTC?��616<�/��g HS|?z��as�������1��?��0�?c�r AW$O��!`��%rzP<]O��t\awxOV4 �`�O�$�a�O�ҵ��O`����O��.EN _p�D�`<_��ite_?���v t_�� aO��IF{?�Ԉ`����) "s_�Ep�a�O-�>n1!Ot�.vTo5!�_��F8���o^837�o*QogW-���o�/��X@�PDT4��_&��ze�OHf4�_\79���MN������f�tro9?6�rx�i0���J59L��%����Ak��P��&��_p�o�Fp_-o`�@�?(�f1'?�pm_d��O0��ٟ�O.�pe����m\�A��/_���N��2.p�͆cW_��֮͠c�a/\ �R8���(Las $���O_���0x���bo��<����I�̿�"% ���K��/?�s�if<Ϟd�?�NT+���Se����/�/�C/�����'37̏�iUf\����$S<G��Ԁ6h��RD�YLS߱�oI�om8w��_#�ps0������hVmj��93����E�ogW�P��ch\?�I��ퟓ�q �o����rvi7߂]S�/������V(s�t,��F���@�t	l�u&5/�����T
�hWi��ݶSe0��6O��sr��	�&�! ��y8P`��dr׏�o3PR	I���a�O�/	9X/��spr�ߕ�����Li?/��3 3H6x/�d94'��963�q54 H�/vg653�/r4 H���&0�/�'��� X?�v72�Ie?�g1I3;?��7�/58r?2�'6�/��Lo�_��t �ͅA�ϐOc�m�osK�!����O�����,�O9��O�OS�ualP_��8�?a_?�g8�_��wr+��j83�?!�_]�&��NDSO-�f7O=��!�Y�ad�O9k1l�o�s_#1�o���ip#�-Et�op�RI�N,��/I���V�A�=SE_��0�
S���Z 0+ͅcmg�Z��0 4@�"�ut[/�of��`�M�r����@�����596O_��4DЏ��U��#o(� I�c5%r_����e`���G�������c���AL"���lga33_U�oy� -<�t
��	e�@t���RTU���h�z�xo��vo;��'O�52 ����4��'�2Yu\�� vOA���42I`FĿ
d -�ݕE��� (o�[��"E3�yo��Wel�_��������WMG��Ϣ3aP@�Ϣ3wm�g[����߂�- ����On�45�?�fCqMk�IO��  �� �������1���2�g��y� R�;�Co���4(S�`�⯔��Ġ��3IF���� 1!(�z�0at��cNT��q���R8�Ϙi5᯳W2\��� O��W?��˿ݿ�0���7��4SiZ/<�0�=�K�!�cl�i5c\sw/�S�AD�f��CVt�Dt.�Q�mt�_�e���V��-V�  /6��Nlo���1��\�O�/C@ �/�4 �/�i�0e/�/1_�W62˟���o�/�eJ7��esrv�?�) "�?�svh�?
o�N� ��?�.p[�tvh9moO�U749LORp`r��OutlO?�t\�?��j�_�/x/�/h_ mpc��&y�9\KO�j�_�/��_�uXP�/D�H18gO}�oOnn�O�%N�߬u�'o���n]`8���oRCM�o�u�n�_��$./_�#��m  �H552�ab�e�q38BSR�78�p�q�r0��l�ibJ614~�cATUP�@wrmc�p545zP�sgt�r6��VCAM�3C�RI�p\rc�pCGUIF�  �q2�p�td.f�NRE�N rco�p631�  - Pr�pS�CHV� DioDOCV>aIFL�WCSUJ18�0�p�1}�EIOCk  ��4�p54�p�R�`4�9�pgm�S;ETf�Sta�q�q/lay,�p7�q�0MASK�S�PRXYZaa�p�7f�C�pHOCOC��3.3�r�p\c΂51�p��qoapp.�q39f��j50�q�ust�3�LCH��A`
OPLG�1"�E��� "L3�MHCR  08 (Ā�S@�Reg��CS@�p�1H��p��q5�p�08\�pMDSW�  URGw�MD����sOP��\!�MPR�ra�4�Հ!��o�f��p! p��PcCM�H��R0БPath���p@aH�"ՀRm����pTP���nՀ816�50�p�g��āS��ol,r�9Ղ:�FRD�p�(Q�pMCN��cc��H93�pLNP���SNBA@�rSgHLB��֑SMx�7lrn?�63�p�r�q2�pL�HTC�pX�TMILVs�r�LT��PAu�Y�sȡ�TX>aEN��ELU�th��0�@`��8�qHѰr9��`ρ9�5�p �Հ7��U{EV��adin(�qC�����pUFRI�;eeO�VCC�pt��VCOY���VIPN��spd�[�I^��p�X͡tsπWEqB�p��?�HTT�p� L2�R62�pC�oo?�CG��d��IGt�
PRIn��PGSN ng�wIRC��ne ���H84�prd6�R�7��@�R��L�53^�p\lcl�q8�p�D" #4�6M� ���52�8�R65�9��|�5�r d K�6��p��4�49�Yp`S��p5�̰L�06�p�VG MD�o�g,� ��66�p��ðA{WS�pJ643��LIက�V��pzdҡ��u�GD����q�,%�h�TY�� ����TO�p<q�q6�g��|� �-@��ORS\Y��R68�p3��sOLp�ģOPIɰ�sguK�SENDH�/аpLP�T�S��\y��ETSɰ2!��6�U����-�43� !D�VRu�ryn:�IPN��onF��Gene��oaytD (S��E��ցI�0�֙���p�yttw\sg��g "�֏�6h��L�yt\str�ոA�ՀA��hk_t���yt�����es�լr��j7��mon.�՜A��
d@6��s-@�ׂ�yt�46\�`Q���qh83��zDlli4�F�clc�`�$rt{� ���¥���yt��w�x��U�Ӑh8��nde���AxV絰����N���ͰH��epen���yt�T��Ģ���ob3攢��h89Ԙ���p��Pv�ed�����4 J7R8�05��0l��ձ`"�t644����� #II���r�p���Ճ"S��/л%��5;94G�tom���!�R J��� 6��Se3�ar3�E��t32�%�QsysG�F ��������wetr��urnk�����20�x78���'�rn6����6�\jtET��
;jo��ta.C����gr������� ����<���ge���017��2�yt�yt75b���Lj(���]7 "P��T`dc��) ��	�`���r��1%at�b@O���p��daW(?�4tv/ 4oh��c�8}���s?yR�?�=l�ogm�?�;ild�?1<d�?N�@���H0@O�M���p1|O��;x@���ytV��1����O_�	8�aicC 2�9����C��7��6�E �� `E?k3edg?y=wm�`O�Rhl$_�2G&heh>�m_��7�5l�O2 24O Oaw4OJmsdh\o�;dh2����osqz�o�kl@���o�o��:��+F�cet�'-�6J8"W<Q��1 (F���pbDa�0��fr{F�� �� �f22.fv�FusS�pkg�M!INgD�x����,��u��o�{��5s22�xsiRC��n VM��^�99�2�W� ��J9�b��st�'T��O 92\�6CMR/d#Z��O;��ݎv'���t�mF����f8�va%t��t+9>e��6ft"/��z_v(��ɟ?�4o���,���կK����vs�w�8��Dni�o��lb��蟮���p��W�\���vsmTڴaz�"����οD��of���ow�L(ώ�slw���f����e�w�����*�vrh�ys�+N3GeN��v�Y25:�oad��(Na�NJ?��nd�� "NwV w �(F8����rrd�6`��lAe&���C�U�4;���Ok7\��8���rk&,��gl��P��1g�Gt��il��������  � P2^���38��rC ����0��J614��ATUPj���5�45����6F��VCAM��C�RI!7� , UI�FB���2��ans���CNRE�'��6�31��RI��SC�H�u65DO�CVN�ns� CS�U�T|���0��HA�EIOC% "v��54��R69�65\� ESET��W�����7 {Cu� MASK��t 1PRX%YUJ N 7�ל�OCO�om�513r�,,������ ��98\t����]��[39�v!��o�ftwLCHz!g�OPLG:�-950ai�P\]P��e f,S�r��CS���^g_lo��5�� �pDSW6�rs70<!Pl DKcOPP4�PRQGS01� n Ad�����X#PCMAa� ��0�%���v�dv; �A
T�X��0��1AD#IG� �!H ,�S�r723��98AU�+ FRD!h#�RMCNr	H93z��R2SNBA"��C+ SHLB�	S�Mp5�n m�J;52�HTC���oTMIL6�Se���PO�0PA�8�6*TPTX�VR��0ELA4ool,���� P��8��\�sv���qSRV�T��95Q$95�A\et� UEV��@a\AC!]�[AF�R!r��C!o;l.�VCO��P.��VIP�4e�� mI�t34[SX�>��WEB���@E(�1T��,�l2ttQ, G�Eg\tk�IG�E#@`PPG�S"�PRC�4"T�AN��84��#R-7�taQR�(
�R53�tRJ698��R66a�52a- E��R{65qr Im��5a��l��573R64q���q�5`M� 061%�BF�f�R   ���WS!40�AC�LIQf9�PSniKaMS�E�Rn`n��597{1TY�4o76 J, TO��tL���6�9 (k�5Pfer@OR�S�CR68��\�sn[!L%CSN� OPI1Tp�\0� ���sn.��L�E ��bS�fX�0ETS 1T����h#�0a�P. FVR� �,Q�N�4�GeneN�a
@�D�x���yMG" �y���y�g_cc�y"�xc�mg_�y��yvth�yR�x3(�,�>��P�b��z1��z! c=v�yon T�yh" �xhr�x�b݉1�`]��iA�y CV�yCP �z��x��xt���	q�ypse������wr57� In����xy͉576��(�p+�)� ����L� �"Al��w6\ab,����j8<�B��lh ��PR<�J8�z�PxC;�8�J�psr��P��x96\{� (P�y�����A�xY`�� -��iv{�R �DM<�H7�zH6�{66�3�1�x�[�tor������(�y�m�!��sZ�r]�2����nalۺ2��)�޸stK��}gstr��ypsk���=�\p����xj932|�C��}�)�x8R�x2}����ʙ.|�޸_w���}hk_k�FH��z9!�xkke*�n�95
����yhe�z885,�f�l.��H��et_w�y�"M�c0� �� �zbak�H��Z�ent��h�\m���s���� ��d �༛�Y�;�(�Z�@�z9Pf�yv�@��.� ����� l�n�( l�gd��=
i��!� Z���+�00iB\�H[�H���� -ڽh[�C" #��8e2��2�@}�OR��8� ���iB/̿N&@�"F���f��h@�+�=���tk� OR�����83�i1�t� ˚�~nc+��f�c����5���83A5�z����i�;�5:l�B�ri��ER���b݉ (ˊng,(�@�,4�*RȭY�k�xmo�`]/��9p�+��ptp�z(��5\pk�=O?�A�45[ڈ��0�/�/ ?S�i�k߽�ij��
���?�+�db��� s50l�a��x���S�[d G�yϋ�cce��0K�50�Kz1�y�6h�Je�RDE��yqI;nt�
 Pa��(��9\g{�H�919p[�p�\:� Vi��tool<?ވ	�J�[�uppK/=_��vk{��K[��Z��Z� �O�O�O�8�OK�H��?ξ�_rj;*h�nd9r{�H]end��I�r:�(�3��o>�7!3;���/�&7;*� �{X�j�|���"�4�?  am_xO�#ve�ʘ���vI����o�?|�xj{��� r�Tz{�] R5;�;J9�;989ﭹP���_��p�m
�
�`�����e�kR Rl�}++R7�J L:;�) "���Kz�/p+zx�d	�-�|�	��633�06 Sl�I~R6�st�z���:�LND��IF� K�45��-co�n{
C9�i�*ar� �jyp�	�ds �"����ENl�y���s��l�gr��e9-����856��`��zrpi{�x=H�4� l�^�wj�!� r˛vv�:nn��}RC:| �� �J9�Z����867�13J;6��8 �J�T�`��(iR��R�|"ٟc  �STD��.p?LANG&���
��r��ti����P��hq��)0-�� E��Okg
��y` ��y5����R730���(��8 (i��E�rrP��,�`��P�C��x���rvge`������8���ge���a<����	�.��i�sio��ckin�� �R�(���pGi� �����؁��yj	��PFK"���XA��\@��BP4���!��d��aabbPbbb�����P`��P��(1��SP��Р�FS J��J�91��6859X!	��02*4<627���Y���,����X���s\�GFSO������sex��/�v�r�����&���R]G(R68'6�4����#8	G =(� CCR��I����cc�� "C�kH���9�\R�BT}rgOPTN�4�4�2�4�?x�?O"Ocrg.8E�F��8E��
D�PN��d�uDio{n tEnd.tE�xa�FINTtE��7tE� ntEa�@tE�0�"tEHQtEhd\mƘFHD�F�uD\eCrh�F���O�AitEp��sF�"UiretE0huDtuDrh�GdCted �����򭔏n An�U�Y9p9 �Ut2��8��0E���a�U�`t f�1���2��� m�U�a�U葠U�-`s�U�ѠW
 ��1�����6h�U wR88�U851_fy4�`�Utiar�U���it� ��l"���MR S�f`�fTcXP�U��epm�f�" #1�f! T�fy��fm�g��e�P��U 2�U 70�Uo�njg���@_f J�7�Vipp�fon,��U���X�v4��j7�9�fc��e]h98xjg�"��\chp�W�EN�vd@Pb{St�o'�� E f�@�VgF0�el�gxѠU���j8svY��f���6�uharel�UKA�Ro�Comc�u�R�ĆL*wp\ �V
t+vY�u�fp\e�V�AN"���k�gpcp_f1a!I�[�f�4y�wf
! Gf ;Co�uarwf��FІ84_f5 H�fH84�v63 �H�fH7�v779�_f24��7rw69V*�65�f1�g8p�v�V75�VIC �fw AP7v893�`��R0���B�eck���Hs�
E����#fMNS+v�ПVՐ�V�P_f-]�_�Q�V8X�\���tch믅��U3\pSfWT"p_fdBe��Zhin_�� �03jgoX��(7ROB�wOG���A�Ue�A�^�HR�Px`flRuuyQuug_Sfz̉3uh523.�{le*writy ��6�2�6�5sv554f�4І40����H60�v0�h�[�08��+�=�O�a�b��8< ���68v�`��s�75^0��A�rw7��h����וл��3�v3Y� &� �େ2f���� 29#f�p����\ib<f��;sbs8�w��o scbP1o�Cja��Ly2%� -k�E"�74�9 wf� (W_�	`��XPLF���wvF�E�X�φ�`we�Vp��a\cwvTf͸�z50+�G"WV����֤u���2�Y �� ��nte�g�����f04 (��gx��D����BP	Xk���I/��`o�!d�@��G��pv �kϥ�ib�hp 
om �wfE�A�f��&Hfdn���z8Z�0f��ؿ�ra�W�_��oi �<�al�VV�Ax�V�2�� 996#fVCA��,�vast#/�q� ��"��dp/fyn:�f�i���58����D��odif��.e8�DP��q (d��o "���o��Rg�d98Ԑ'G��strS����OAW���wR73��v16"� Rf�7�9�2���iTra���c�h�/�wv"�TP+v̀��tpe��c�wor���+R�C�59�8�� S�5+�809�?��C��f�"z\mߦ<�����RE��$sFL&0�pcz��6�verv�gng�_��746�_��S�_� Ch�?�� ����8th\��0�897i3�g]���6�f!��by$�x���� T��w��&w& ���rk����`s�H��VAGǧset�99�������$FEAT_A�DD ?	�����q�p��	 x������*� <�N�`�r��������� ̏ޏ����&�8�J� \�n���������ȟڟ ����"�4�F�X�j� |�������į֯��� ��0�B�T�f�x��� ������ҿ����� ,�>�P�b�tφϘϪ� ����������(�:� L�^�p߂ߔߦ߸��� ���� ��$�6�H�Z� l�~���������� ��� �2�D�V�h�z� ��������������
 .@Rdv�� �����* <N`r���� ���//&/8/J/ \/n/�/�/�/�/�/�/ �/�/?"?4?F?X?j?�|?�?�?�tDEMO� ^�y   x�=�?�?OO %OROIO[O�OO�O�O �O�O�O�O__!_N_ E_W_�_{_�_�_�_�_ �_�_oooJoAoSo �owo�o�o�o�o�o�o F=O|s �������� �B�9�K�x�o����� ��ҏɏۏ����>� 5�G�t�k�}�����Ο şן����:�1�C� p�g�y�����ʯ��ӯ  ���	�6�-�?�l�c� u�����ƿ��Ͽ��� �2�)�;�h�_�qϋ� ���Ϲ��������.� %�7�d�[�m߇ߑ߾� ����������*�!�3� `�W�i������� ������&��/�\�S� e�������������� ��"+XOa{ ������� 'TK]w�� �����//#/ P/G/Y/s/}/�/�/�/ �/�/�/???L?C? U?o?y?�?�?�?�?�? �?O	OOHO?OQOkO uO�O�O�O�O�O�O_ __D_;_M_g_q_�_ �_�_�_�_�_
ooo @o7oIocomo�o�o�o �o�o�o�o<3 E_i����� ����8�/�A�[� e�������ȏ��я�� ���4�+�=�W�a��� ����ğ��͟���� 0�'�9�S�]������� ����ɯ�����,�#� 5�O�Y���}������� ſ����(��1�K� Uς�yϋϸϯ����� ����$��-�G�Q�~� u߇ߴ߽߫�������  ��)�C�M�z�q�� ������������ %�?�I�v�m������ ��������!; Eri{���� ��7An ew������ ///3/=/j/a/s/ �/�/�/�/�/�/?? ?/?9?f?]?o?�?�? �?�?�?�?O�?O+O 5ObOYOkO�O�O�O�O �O�O_�O_'_1_^_ U_g_�_�_�_�_�_�_  o�_	o#o-oZoQoco �o�o�o�o�o�o�o�o )VM_�� �������� %�R�I�[�������� ��Ǐ�����!�N� E�W���{�������ß ������J�A�S� ��w����������� ����F�=�O�|�s� ���������߿�� �B�9�K�x�oρϮ� �Ϸ���������>� 5�G�t�k�}ߪߡ߳� ��������:�1�C� p�g�y�������� ����	�6�-�?�l�c� u��������������� 2);h_q� ������. %7d[m��� �����*/!/3/ `/W/i/�/�/�/�/�/ �/�/�/&??/?\?S? e?�?�?�?�?�?�?�? �?"OO+OXOOOaO�O �O�O�O�O�O�O�O_ _'_T_K_]_�_�_�_ �_�_�_�_�_oo#o PoGoYo�o}o�o�o�o �o�o�oLC U�y����� ��	��H�?�Q�~� u���������׏�� ��D�;�M�z�q��� ������ӟݟ
��� @�7�I�v�m������ ��ϯٯ����<�3��E�r�i�{�����˽  ¸��� �)�;�M�_�qσϕ� �Ϲ���������%� 7�I�[�m�ߑߣߵ� ���������!�3�E� W�i�{�������� ������/�A�S�e� w��������������� +=Oas� ������ '9K]o��� �����/#/5/ G/Y/k/}/�/�/�/�/ �/�/�/??1?C?U? g?y?�?�?�?�?�?�? �?	OO-O?OQOcOuO �O�O�O�O�O�O�O_ _)_;_M___q_�_�_ �_�_�_�_�_oo%o 7oIo[omoo�o�o�o �o�o�o�o!3E Wi{����� ����/�A�S�e� w���������я��� ��+�=�O�a�s��� ������͟ߟ��� '�9�K�]�o������� ��ɯۯ����#�5� G�Y�k�}�������ſ ׿�����1�C�U� g�yϋϝϯ������� ��	��-�?�Q�c�u� �ߙ߽߫�������� �)�;�M�_�q��� �����������%� 7�I�[�m�������� ��������!3E Wi{����� ��/ASe w������� //+/=/O/a/s/�/ �/�/�/�/�/�/?? '?9?K?]?o?�?�?�?|�?�9  �8 �1�?�?	OO-O?OQO cOuO�O�O�O�O�O�O �O__)_;_M___q_ �_�_�_�_�_�_�_o o%o7oIo[omoo�o �o�o�o�o�o�o! 3EWi{��� ������/�A� S�e�w���������я �����+�=�O�a� s���������͟ߟ� ��'�9�K�]�o��� ������ɯۯ���� #�5�G�Y�k�}����� ��ſ׿�����1� C�U�g�yϋϝϯ��� ������	��-�?�Q� c�u߇ߙ߽߫����� ����)�;�M�_�q� ������������ �%�7�I�[�m���� ������������! 3EWi{��� ����/A Sew����� ��//+/=/O/a/ s/�/�/�/�/�/�/�/ ??'?9?K?]?o?�? �?�?�?�?�?�?�?O #O5OGOYOkO}O�O�O �O�O�O�O�O__1_ C_U_g_y_�_�_�_�_ �_�_�_	oo-o?oQo couo�o�o�o�o�o�o �o);M_q �������� �%�7�I�[�m���� ����Ǐُ����!� 3�E�W�i�{������� ß՟�����/�A� S�e�w���������ѯ �����+�=�O�a� s���������Ϳ߿� ��'�9�K�]�oρ� �ϥϷ���������� #�5�G�Y�k�}ߏߡ� ������������1� C�U�g�y������ ������	��-�?�Q� c�u������������� ��);M_q ������� %7I[m� ������/!/ 3/E/W/i/{/�/�/�/ �/�/�/�/??/?A? S?e?w?�?�?�?�?�1�0�8�?�?OO 1OCOUOgOyO�O�O�O �O�O�O�O	__-_?_ Q_c_u_�_�_�_�_�_ �_�_oo)o;oMo_o qo�o�o�o�o�o�o�o %7I[m �������� !�3�E�W�i�{����� ��ÏՏ�����/� A�S�e�w��������� џ�����+�=�O� a�s���������ͯ߯ ���'�9�K�]�o� ��������ɿۿ��� �#�5�G�Y�k�}Ϗ� �ϳ����������� 1�C�U�g�yߋߝ߯� ��������	��-�?� Q�c�u������� ������)�;�M�_� q��������������� %7I[m ������� !3EWi{�� �����//// A/S/e/w/�/�/�/�/ �/�/�/??+?=?O? a?s?�?�?�?�?�?�? �?OO'O9OKO]OoO �O�O�O�O�O�O�O�O _#_5_G_Y_k_}_�_ �_�_�_�_�_�_oo 1oCoUogoyo�o�o�o �o�o�o�o	-? Qcu����� ����)�;�M�_� q���������ˏݏ� ��%�7�I�[�m�� ������ǟٟ���� !�3�E�W�i�{����� ��ïկ�����/� A�S�e�w����������ѹ�$FEAT_�DEMOIN  �ִ���ΰ��INDEX������ILECO�MP _���7���-��SETUP2 �`7�A�� � N l�*�_AP2BCK 1a7�?  �)Ҹ��"��%����ΰ:��� ��Ե��*߹�N���[� ��ߨ�7�����m�� ��&�8���\��߀�� !��E���i������ 4���X�j������� ��S���w���B ��f��s�+�O ����>P� t��9�]� ��(/�L/�p/�/ /�/5/�/�/k/ ?�/ $?6?�/Z?�/~??�? �?C?�?g?�?O�?2O �?VOhO�?�OO�O�O QO�OuO
_�O_@_�O d_�O�_�_)_�_M_�_ �_�_o�_<oNo�_ro�o�o%o�o�oF�z�P�~� 2��*.cVR�o�`* �F�cLpZepPC�x��`FR6:D��~\��{T� �'��u�Q����w�Yf*.F
���a	�s��Ռd�����STM �"�-��p��Y��`iPe�ndant Pa'nelY���HO����?���[�����GIF�6�A�"�ߟ񟆯��JPG����A���0c�u�
��zJS�=��`У+��%
J�avaScripti���CSZ���@����k� %Cas�cading S�tyle She�ets�_`
AR�GNAME.DT�lD�\0��P��`�q��`�DISP*g�J�D����σ�����ϡ�	PANE3L1��O�%D�8�x�k�}�+�2m���b� ��~ߐ�%�0�3��W�@b�E����0�4u���b�����-�(�T�PEINS.XML4���:\H����Custom T?oolbar�����PASSWORD���}nFRS:\����� %Pas�sword ConfigXoV�� O��o�?��u 
�.@�d�� )�M�q�/ �</�`/r//�/%/ �/�/[/�//?�/�/ J?�/n?�/g?�?3?�? W?�?�?�?"O�?FOXO �?|OO�O/OAO�OeO �O�O�O0_�OT_�Ox_ �__�_=_�_�_s_o �_,o�_�_bo�_�oo o�oKo�ooo�o :�o^p�o�#� GY�}���H� �l������1�ƏU� ����� ���D�ӏ� z�	���-���ԟc��� ���.���R��v��� ���;�Я_�q���� *���#�`�﯄���� ��I�޿m��ϣ�8� ǿ\������!϶�E� ����{�ߟ�4�F��� j��ώߠ�/���S��� w߉���B���;�x� ��+�����a���� �,���P���t��� ��9���]�����( ��L^������� �$FILE_�DGBCK 1a���� ��� ( �)�
SUMMARY�.DG�hMD�:�0t Di�ag Summa�ry1>

CONSLOG&	t��CConso?le log�=	TPACCN��/%�4/?TP� Account�in�>
FR6�:IPKDMP.'ZIPh/l
�/�/�@P Except�ion�/n+ME?MCHECK*/��@?�Memory DataA?��LN�)	F�TP��?'?�?K7��mment T�BD�?u7 >)�ETHERNE�T�?f�!OHOC�Ethernet� �figura��/D�1DCSVR�F�?�?�?�OQ1%��@ verif�y all�O�M�,��EDIFF��O�O�OO_R0%�HdiffQ_W�!>�@CHGD1F_-_?_�_ f_�_S+P�Y2�_�_�_Xo� �_ooGD�3No5oGo�o �no�fUPDA�TES."pi�FRS:\ a}�DUpdates� ListafP�SRBWLD.C	M�hLr�c��PS_ROBOW�EL�?<�aHADOW�o�o�of�Q3�Shadow Changesi�ޗ�=�&�NO�TI�OA�S��O5NotificqB<���O�AJ?� nc��p���D��L� �󟂟���;�M�ܟ q� �����6�˯Z�� ~���%���I�دm�� ���2�ǿٿh����� !�3�¿W��{�
ψ� ��@���d���ߚ�/� ��S�e��ω�߭߿� N���r����=��� a��߅��&��J��� ������9�K���o� ���"�����X���|� #��G��k} �0��f�� �,U�y�� >�b�	/�-/� Q/c/��//�/:/�/ �/p/?�/)?;?�/_? �/�?�?$?�?H?�?�? ~?O�?7O�?DOmO�? �O O�O�OVO�OzO_�!_�OE_�Oi_{_�$�FILE_LpPR�[p��_P�����XMDONLY 1a�U~ZP 
 �
_ �_._oR_o;o__o �_�o�o$o�oHo�o�o ~o�o7I�om�o � ��V�z� !��E��i�{�
��� .�ÏՏd�������� *�S��w������<� џ`������+���O� a�🅯���8���߯~�ZVISBCK�X|�Q�S*.VD�|0���FR:\���ION\DATA�\�â��Vi�sion VD file\�j����� ̯ڿį�����4�ÿ X��|ώ�ϲ�A��� e�w�ߛ�0�B���f� �ϊ�ߛ���O���s� ���>���b���� ��'��������� ��'�L���p������ 5���Y���}���$�Z�MR2_GRP �1b�[�C4�  B� 	 ��Qk}h E�� �E�  F@ �F�5U�/
h L����M��J�k�K�v�H�,�Hk���?�  �/h 9�tQv8����6h�%�A��  3EBHeB)�a `�E@i/�g��h @UU�U�U��>�]��>П�;r�8	===E���<D�><��ɳ<�Ε�:��b�:/'79��W�9
@�8�8�9���T/�Q/�/eE7� E?p D�D��/�D�  D��  Cζ/9
_C�FG c�[T ��/?0?B?�N�O �Z
F�0x1 }0�RM_�CHKTYP  ��P� �P�P�P���1OM�0_MIN��0
���0�P]X�PSSB�#d�U�Pi�?	��3O$O�UTP_D�EF_OW�P
|�Y?AIRCOM�0�JO�$GENOV_RD_DO�6�RnxLTHR�6 d�E�d}D_ENBiO �}@RAVCGe��7� ��Fn�H E�� Ga� H�� H�?@Jh`�/O�?_�G_X_{ ���AOU�@kN� {NB{8���_y_�_�_�_,� � B�a �%o�? doCOm?aUc~	��Y+O�@SMT�Cl��IZ �0 C���HoOSTC�"1m�o� 	
xM
{
:byeV���� �zu� ��$�GH���p	anonymousK�y������� ��	-�A�c �V�h�z������ ԟ����M�_�@�R� d�v���ˏݏ��� �7��*�<�N�`��� ��������̿�!�3� �&�8�J�\ϟ���ï կ׿��������"� 4�w�X�j�|ߎߠ��� ���������0�s� �ϗϩϫߜ������� �����K�,�>�P�b� ��s��ߪ��������� G�Y�k�L�p�� ������  $6YZ��~�� ��	�-? /S uB/h/z/�/�/��/ �/�/�/
?-/_qR? d?v?�?�?��// ?�?I/*O<ONO`OrO �/�O�O�O�O�OO3? E?&_8_J_\_n_�g�a�ENT 1n�i��  P!�O�_  �@�_�_�_o �_+o�_Ooo[o6o�o �olo�o�o�o�o�o 9�oo2�V� z�����5�� Y��}�@�v�����׏ ��������+��T� y�<���`�����埨� 	�̟ޟ?��c�&����J�QUICC0���p�!172.8.9.225�����1�����3���2�4��"���!ROUTER��`�r�ӿ!PCJOGԿ���!192.�168.0.10�����CAMPRT,$� �!�1�K�2�RT��O�a��ψTNAME !�Z?!ROBO=����S_CFG 1m��Y ��Auto-sta�rted�4FTP�?[��?�O��O �߼������ߋO�(� :�L�o�]����� ������04�F�X�9� l��P���������z� ������#F���Y k}����?�?�? �?.b�CUgy �N����� �-/?/Q/c/u/�/� �� /�/6?)? ;?M?_?"/�?�?�?�? �?�/p?OO%O7OIO [O�/�/�/tO�?�O
? �O�O_!_3_�?W_i_ {_�_�O�_D_�_�_�_ oo/orO�O�Owo�_ �o�O�o�o�o�o�_ +=Oa�o�� ����4oFoXojo K�~�o��������ɏ �����#�5�X�ڏ k�}�������ş�� ,�>�@�1�t�U�g�y� ����`���ӯ���	� ,���?�Q�c�u��������_ERR o��ʡ���PDUSI�Z  3�^L���ȴ>�WRD �?"���  �guest -�!�3�E�W�i�{����SCDMNGRPw 2p"�˰���3��-�K��� 	P01.o05 8�� ������>0�j  �2�1�� � ����T���������������$���ϿQ�<߬u�`�������  �  -
��N(�P,�(�����Q���m������l��- 8�#{�d������"ߙ�_GROU���q������	�����4S�QUPD'  �ȵX��TY�����T�TP_AUTH �1r�� <!iPendan�����8�g�!K?AREL:*����KC-�=�O�%��VISION �SETb����3� #�������"� �� _6H�l~��CTRL s������3���FF�F9E3��F�RS:DEFAU�LTFAN�UC Web Server���� 	�Ĵ}��������WR_CON�FIG t�� ���IDL_�CPU_PC*�3�B��I  BH�/%MIN:,��M%GNR_IO������Ƿ1 NPT_SI�M_DO&�+S�TAL_SCRN�& ��*TPMODNTOL�'�+bRTY�(I!�&����ENB�'��-$O�LNK 1u�� �Q?c?u?�?�?�?�?>52MASTE~ ���52SLAVE �v��34��O_CFG�?IUO��OBCYCLE>OD$_ASG 1w����
 �?�O�O�O �O�O�O__1_C_U_�g_y_�_�;tBNUM��Ĺ
BIPC�H[O��@RTRY_CN*�"ĺB�!(���P1�ȵ B;@Bx�>�Jo�1 �SDT_ISOL�C  ��f��$�J23_DS4��:��`OBPRO�C?�%JOG^�1�y�;��d8��?��[�o�_?؟֟O|QNs��@V����-�~o��h�`Y A�_�bPO�SRE�o�&KANJI_�0���/k�+�?MON zg��2�y�Ϗ����HҾ)�0c{,�9�<T�f�CL_LY �R��_k�EYLOGG+IN@����ȵ��$LANGU�AGE k2e$ 㑱�LG1bY|�2���3�x�ʗ���O � '�0,�� �
q��3�MC:\�RSCH\00\���LN_DISOP }�?f�M�Km�OC�"@"Dz�h#�A�OGBOOK ~K��w�0��w�w���X��� -�?�Q�c�u���11����	���h��޿����ॐ_BU�FF 1@= ���)�����E� a�sϠϗϩ������� ���B�9�K�]�o���ߓߥ��ߜ��DC�S �� =��͗�ֿM�l:�L��^�p���IO 1��K No�� � �����������%� 9�I�[�m��������� ��������!3E�Y��Ex TMlnd ������ 0BTfx��� ����//����SEV`}��TYPln��/�/�/)-P�RS�P���b�FL 1���`��?,?>?P?b?t?��?�/TP��loq">��NGNAM�d���Ւ��UPSu�GI��U\�e�1_LO{AD�`G %}��%DF@GI6��?�[MAXUAL�RM�Wk�X\@�1_PR�T`ԣ��Z@Cx��ꩦ��OV�x9ŜC�`P 2��K� �9�	q!>P]  ��OQ� R9_$_6_o_�]_�_ �_�_�_�_�_�_oo @oRo5ovoao�o}o�o �o�o�o�o*N 9rUg���� ���&��J�-�?� ��k�����ȏڏ���� �"���X�C�|�g� ������֟����ݟ� 0��T�?�x���m��� ��ү��ǯ��,���P�b�E���q���SGD�_LDXDISA��0�;��MEMO_{AP�0E ?�;
 j ���π*�<�N�`�rτ�Z@I�SC 1��; �����T�A���ϛ��$��Hߙ�C_MS�TR �B-g�S_CD 1����<� ��8���������"�� �X�C�|�g����� ���������	�B�-� f�Q���u��������� ����,<bM �q������ �(L7p[� �����/� 6/!/Z/E/W/�/{/�/ �/�/�/�/�/?2?? V?A?z?e?�?�?�?X��MKCFG ��vݽO�CLTARMU_�2��G�B P��2�@>OFD{@MET�PU�C�@��~�N}D�@ADCOL`E��@kNCMNT�O 9tEo� �v��N�5C.A�O�DtEPOS�CF�G�NPRP�M�OYST@1�ޯ� 4@��<#�
oQ�1oU_�Wk_ �_�_�_�_�_�_o�_ oOo1oCo�ogoyo�o��o�o�o�atASIN�G_CHK  ~�O$MODAQC��?���>+uDEV� 	��	MC}:_|HSIZEѽ����+uTASK �%��%$123456789 ���u)wTRIG 1���l#E%��)���`�S�6�%C�vYP�q�>�At*sEM_I�NF 1�#G� `)AT&FV0E0`��׍)��E0V1�&A3&B1&D�2&S0&C1S�0=ƍ)ATZ׏+��H/�W��K���A����j�ӟ����	� ��.���� ���;����Я⯕� ���*�<�#�`��%� ��I�[�m�޿鯣�� K�8����n�)ϒ�y� ����{��ϟ���ÿտ F���jߡ�{ߠ�S��� ������������T� ��+ߜ��a���	� ����,���P�7�t� ��9��]�o��� ��(:q�^��=�����XNIT�OR�@G ?s{ �  	EXESC1�32%3%E4%5%�p'7%8%9�3 �� $�0�<�H� T�`�l�x�T��2�2�2�U2�2�2�2�U2�2�2�3��3�30+qR_G�RP_SV 1� (�a���:��hK=�&�7��);���=>�T�Eav�q_�D{�~�1PL_N�AME !#E�0�!Defa�ult Pers�onality �(from FD�) �4RR2�! �1�L68L�@�1P
d d �?v?�?�?�?�?�?�? �?OO*O<ONO`OrO��O�O�O�O�O�OJx2 e?_ _2_D_V_h_z_�_�_�_r<�O�_�_ �_o"o4oFoXojo|o��o�o�i�V�_�n
�o�oNtP�o*<N `r������ ���&�8�n� ��������ȏڏ��� �"�4�F�X�j�|�K� ]���ğ֟����� 0�B�T�f�x����������Ү FnH� F�� G=�<�'�   �����"d���0�B�&�d� r��׭Ҫ\�������ݿ� ͸���  ��0�6�T�vϿ ��ϩ�ͰA�   ��˿��Ǹ]0���ƿ 3�¿W�B�{ߍ�x߱�dB5K3�9^0`�!0 � ��0�� @D�  &��?����?� ��!A�����$���(;�	l�	 ���p�V� ]0M� � _� � �l�r��� K(��K(��K ��J�n��J�^J&Ǔ�2������� �@Y�,@Cz?@I�@���������N�����f���_�I_���SѬ�Ä���  <��% ß3������!?s8y�
�/�!��x����T� ܌�������}���    �������  ���������	'� � 0�I� �  ������:�È~TÈ=���l��	�(|�����ш����ψ��N@0�  '� ����@2��@����@!����@)���C@0C��\C�I�CM�CQ�� ���ģ�%%����� ��B���@0��lc@� ��!Dz�߀�V�//+/Q/��?�� �H@q)lq�%  ��+���� p�!?�faf���/�/V/ ���/;��8� !?/:� ��D4�� \6Pf8�)0c�\�\��?Lv �$���;�Cd;�p�f<߈<���.<p��<�?�L:��ݧA���d�����?fff?��?&@��@��� B�N�@T��,E�	��	A��� dO�O�7H��/�O�O �O�O _�O$__H_Z_0E_~_�MEF�m_ �_i_�_UO�_yI�_2o��XC��E��"Gd G;ML!o�o mo�o�o�o�o�o�o�o $H��iww9� �_�o�U��*�<�ڪ����/�6���@���ď��菎�A�!A�����C؏=�ԏ��X��񨑟,�|����  �P��"�@�<��E� C ���s��x�؄�(������/�B�/B�"�}A��#A���9@�dZ?�vȴ,��~���<)�+� �=�G��j����q���
AC
�=C���������� ��p��Cc�¥��B=���ff��{,�I����HD-�H�d�@I�^�F8$� D;ޓܪ�̠�Jj��I�G�FP<����QpJnPH��?�I�q�F.� D��Ɵg� R���v��������п 	���-��Q�<�Nχ� rϫϖ��Ϻ������ )��M�8�q�\ߕ߀� �ߤ߶��������7� "�[�F�k��|��� ��������!���W� B�{�f����������� ����A,eP �t����� �+;aL�pЩ����(����33:��1��%��3�V��/"��(/:/�!4M��T/f/F1�=���/�/4Ue'��T9�-�)�/�/?�/(4?"<]�P�2Pf>�q��?��?�?�?�?�9���(�?�?/O`O?OeOPO�QB�hO zO�O�O�O�O�O�?t0.__R_@[/X_b_��_�_�_�_�_�Q{f �_�_o
o@o.odorj�  2 FnHn"�F��"�G=��1B# ��C9)��@|�@��o �q�o{�E�� F��`�H C�����oA�`��kE�0wGa �O����{?ސ�q* �\d  zqu `�
 � !�3�E�W�i�{����� ��ÏՏ�������q� ��P+�~Y���$MSKCFM�AP  �%� ^f�q�q�p�D�ONREL  X5[��0D�EXCFENB��q
Y����FNC�����JOGOVLI�M��d����dD�K�EY�����_�PAN����D�R�UN���>�SFSPDTYw0�������SIGN����TO1MOT럜�D��_CE_GRP [1��%[�\�O ��O�&��d�Q�� u�,�j���b�Ͽ��Ŀ ϼ�)�;��_�σ� ��LϹ�pϲ��Ϧ�� %��I� �m��fߣ��OvD�QZ_EDI�T��U��TCOM_CFG 1�Q������"�
��_/ARC_��X5ؙ�T_MN_MOD�E��縙UAP�_CPLF４NO�CHECK ?Q� W5�H�� ��������'�9�K� ]�o�����������v��NO_WAIT_�L���׾�NT���Q��{_ER�Rȡ2�Q��1� A��t���H*�P����`�OI�Px ����!8�?0|4��pBPARAM:J�Q���	���7so� =�`3�45678901 �/ *�?/Q/-/]/��/�/u/�/�/�+�7��?<�7?��UM_RSPACEN��'2$�p?z4�$OD�RDSPE㌦��O�FFSET_CAqR�Ќ�6DIS�?��2PEN_FIL�E�0�$��֌1PT?ION_IO
�=��@M_PRG %\:%$*IO[N�3WORK �Χ=�� ���F7�:�Bh�� ��d�@9(7�A	 ��x�A�5��c��0RG_DSBL  \5☓�|_�1RIE�NTTO��9�C��pZ��a�0UT__SIM_DGX��+��0V�0LCT ��%�ҟDx=gT_�PEXh��?�TRA-Th� d���T�0�UP �u^��Ӡ�oo�_:oHi��$�2ǣ�L6�8L@�_S
d d'?�o�o�o�o �o�o�o1CU gy�������I2~o'�9�K�]��o���������ɏ9�< ����)�;�M�_� q���������H�j3@�H1`��XRP� C�U�g�y��������� ӯ���	��-�?�Q�  �2���������Ͽ� ���)�;�M�_�q� �ϕ�d�v�������� �%�7�I�[�m�ߑ߀�ߵ�����X�ϡ!��*��S�H�Z� ?�}������&?������������ +�I�O�m����?@��|��� A�  �� ��������M8 q\����z��d`O�P1� k߀ ��sd`�R0 ��D$@? @D�  DtD?QD	���U�  ;�	�l1	 ��p�s& ' �j � � � �ʉ�� H<z�H<W�H3k�7G�CG���G9|+c	�H
�X�� CC9P/9P�49S;Q9/��9�  ��  1!�}H7 3����/�1/C/�BY�����XQ�^�H�<Pq/ ܩ/�"2��#�3�.�  �  �0��� �  0��6�/?�	'� �� M2I� ?�  ���
=���q?�;�#&�(�3�/��A�?4;"�B�?�NEPO�  'VP3D�b C�EPC��\Cf C�j Cn/@OROߑ  �����D%�%��� �B���FEP�EF˜@XP�E5z��_s/8_#_H_n_�"?�� �H]2�Yl�A�U  �C�H�A�0p�Q?�faf���_�_s_ ��o(k�18�0>oLj- �!adTW�0yfP�h�Y0�yy�3?L�0�T��!;�Cd;�p�f<߈<���.<p��<�?�ij��WA�Eل1d��31��?fff?��@?&+pVT@���=r�N�@T��IuՉ��&q-�0! ��we o�� ����A�,�e�w� b�������я����l����O��CE����2Gd G;�|>�����ß��� ҟ����A�,�e� ����V����د6���@r�#�5�G�Y��Z�  �_�f�������̿��A @A�@%����5�C��Z���/i�?�؈Ϗ��ϳ�UG�P��2]!YNE� CU%�̣��q�����E�@I�!�t�B�/B"��}A��#A���9@�dZ?v���+~��~���<)�+� =��G�(߇Ԁ�q����
AC
=C�����녡�� ��p�C�c�¥�B=����ff��{��I���H�D-�H�d@I��^�F8$ D�;���ڭ̠Jj���I�G��FP<��Q�pJnPH�?��I�q�F.� D��E�τ�o�� ����������&�� J�5�n�Y�k������� �������� F1 jU�y���� ��0T?x c������� //>/)/;/t/_/�/ �/�/�/�/�/�/?? :?%?^?I?�?m?�?�? �?�?�? O�?$OOHO 3OXO~OiO�O�O�O�O��O��(}���3:��O�a��)U�E3��V�_+_9R�xE_W_t�4M��q_<�_t��=ӝ_�_�4Ue'��T9 �]�Y	o�_-ooQo?lJz�P�bP�n������o�O�o�o�o�i���(L7\�mt�B���� �����o��K�9�o�]�/u������0ŏ�ُ�{f���9�'�]�K�����  �2 FnH��F[�Щ�G=��B@P�!�.�C9F��p��@�2���	��C�E��� F����H CA���S�b����@������¯ԯ��?��T��y�C�C��|�C�}�
  ۯ>�P�b�t������� ��ο����(ϧ��� ��m[�~Y���$PARAM�_MENU ?��U� � DEFP�ULSE4�	W�AITTMOUTތ�RCV�� �SHELL_W�RK.$CUR_oSTYL�����OPT���PTB�����C��R_DECSN��teG�A�S� eߎ߉ߛ߭������߀����+�=�f�a�S�SREL_ID � �U�a�u�US�E_PROG �%p�%b���v�CC�R����ax���_H�OST !p�!�����T�`��8�����:�t���_TGIME����a�?GDEBUG��p��v�GINP_FLgMSK����TR�����PGA�� ���{�CH����TY+PEm�y�a�[� ������ !JEWi��� �����"//// A/j/e/w/�/�/�/�/��/�/�/??B?��W�ORD ?	p�
? 	RS��	�/PNSu��~2sJO�
�TE[��?COLu>8�?Z>L�� �P��p����TRACEC�TL 1��U.z� �`��)O|3BFDT Q��U�^@#@D � sckO}O�O�O �O�O�O�O�O__1_ C_U_g_y_�_�_�_�_ �_�_�_	oo-o?oQo couo�o�o�o�o�o�o �o);M_q �������� �%�7�I�[�m���� ����Ǐُ����!� 3�E�W�i�{������� ß՟�����/�A� S�e�w�����gO��ǯ ٯ����!�3�E�W� i�{�������ÿտ� ����/�A�S�e�w� �ϛϭϿ�������� �+�=�O�a�s߅ߗ� �߻���������'� 9�K�]�o����� ���������#�5�G� Y�k�}����������� ����1CUg y�������� 	-?Qcu� ������// )/;/M/_/q/�/�/�/ �/�/�/�/??%?7? I?[?m??�?�?�?�? �?�?�?O!O3OEOWO iO{O�O�O�O�O�O�O �O__/_A_S_e_w_ �_�_�_�_�_�_�_o o+o=oOoaoso�o�o �o�o�o�o�o� 9K]o���� �����#�5�G� Y�k�}�������ŏ׏ �����1�C�U�g� y���������ӟ��� 	��-�?�Q�c�u��� ������ϯ���� )�;�M�_�q������� ��˿ݿ���%�7� I�[�m�ϑϣϵ��� �������!�3�E�W��a��$PGTRA�CELEN  �b�  ���a��w�_UP �����љ�В�  ��w�_�CFG ������a������������׉���DEFSPD ����`щ��w�IN~��TRL ������8�F�PE_C�ONFI�Ш��O������WLID�ө��	��LLB 1���� t�?B�  B4��� ��� ����� 88�?�0�K�0�G�i�k�}� ������������5Ak��� ��2��	�?~��GRP 1����lb�A�  ��333a�A���D�@ D�� �D@ A@�Ta�d+������� 	='����#´#��B 9!�///O/9/s/
?��?����/�/��.�/ =o=	7L�/?�/?P? ;?t?_?�/�?�??�?<�?�?  DzC Oa�
OHO�?XO~OiO �O�O�O�O�O�O_�O�_D_/_h_S_�_�Z!�a�
V7.10�beta1�� �Ax���R�y�y�Q?���Qo>�\)�QB0����PA��SBp���QA�9Sy�b
a�S �_2oDoVoho��Ap���"���o�o�o�o�ة�KNO?W_M  ��־��SV ������5O8J \u_�k}��ҴJ��M]�z�Д�R�	��%%�"��|����# ��u��P@�a��]�a�q�m��Ц�MR]��}��&%O�P�$�ӏ�KST]1 {1���
 4�� vi�Q:��"�4�F�w� j�|�������ğ	�� ��?��0�u�T�f�����������ү��2r� �a��<K��^35�G�Y�k��A4���������5ۿ�����6.�@�R�d��7�ϓϥϷ���8������
��MA/D  ���)�OVLD  ���G�PARNUM  ������_T_SCHy� ���
�����0�UP�D��������_C�MP_�p|�pp'��e��ER_CHK�����j���Ư�RS��oW_M�O{���_���__RES_G���  o������������� ��2%VIz m`�R�4�\�l�� Q������S�ڰ� S�-�9X]S� ��x��S�������S�&��//S�V� 1���a�q@�c?\�THR_�INR��~��r�edމ&MASS�/ Z�'MN�/�#MON�_QUEUE ����f"��a��N���U��N�&��0E�ND1;�79EXEF?75\�BEE0'?3OPTIO$7D�0�PROGRAM %�*%0T/��~2TASK_I{���>OCFG ���/���?"@DATA��s�+K��"�2 ��O�O�O�O�O�O�O _!_3_E_�Oi_{_�_��_ROINFO�s�oM�
4[_�_
oo.o @oRodovo�o�o�o�o �o�o�o*<Nh`�W�T�oL �	l!A�K_%A�+I�^�vENB|б}����v2��xG%A2�~�{ P(O�4�F� C�e��z�_EDIT ��+O����DWERF�Lg8|# �RGADoJ ��:A����?"���!߆1�q��]��?����A<@��v%�<�l�ӈ���q2��)��R	H0le�|{"6�?
��AF$w�t$ܖ*�=/� **:��"� ����d�1�f�Ցd�[�BU�#���3�E� s�i�{�������߯կ �a���K�A�S�Ϳ w���������9���� #��+ϥ�O�aϏυ� ��߻��������}� '�9�g�]�o��ߓߥ� ������U����?�5� G���k�}����-� ���������C�U� ��y����������� ��q-[Qc� �����I� 3);�_q���t&	>O@/Հ./g/ R$ݙ�/ߓU/�/Q/�/��/�PREF ��)�ՀՀ
߅I�ORITY�72F�>�MPDSP�1я�G7UTFǓކOD�UCT
A�:��/��OG��_TG�΀B���2TOEN�T 1� (�!AF_INE�q0OG!tc�pO6M!ud�%O^N!icmXMOu��2XY"�Í�;�X1)� ��O�OX0��O�O�E�O )__M_4_F_�_j_�_ �_�_�_�_o�_%o7o	*�3"��=Y�yo�o^��>��J��!/�io�o��������AK�,  � 0�q'9K]X5�7��pHANCE !�)��rrn{d�o��uyw	3�?"3ق��PORT_NUM�r3X0���_CARTREPR0|����SKSTAq7� C�LGS @�ȍ��K�X0Unothing� ����̏܌�����#���?k�TEMP �ɕ94����_a_seiban�/ ���/��͟���ܟ�  �9�$�]�H�Z���~� ����ۯƯ����5�  �Y�D�}�h�����ſ ��¿����
�C�.� g�R�wϝψ��Ϭ��� ��	���-��*�c�N� ��r߫ߖ��ߺ���� ��)��M�8�q�\��|6�k�VERSIP0��7�� di�sable�r<�S�AVE ʕ:	�2600H84%4����,�!�.�@�_Od� 	��{2 /����X�e����	�-;
��c�n ��L��_�0 1�
�K�� "��x��0URGE�paB�0T6>5�WF� #DOr6�r�6W�0��"�WRUP_DELAY �;��R_HOT �%%&~1��+R_?NORMALy�2x���SEMI���"/�!QSKIP���w�x��g/�� �/�/�/r-�5�/�'�/ ??(?�/L?:?\?�? �?�?l?�?�?�? OO �?"OHO6OlO~O�OVO �O�O�O�O�O_�O2_  _V_h_z_@_�_�_�_��_�_�_���$RB�TIF?�RCV�TMOUT�B�]�`DCR��E)� �~!7����C���C�?��A7�f�/|#�lD��i���$�a9r/�o�o� ;�Cd;��pf<߈<���.>�]�>Ѓ���o��o'8} 8^p��� ���� ��$�1%�RDIO_TYP�E  �.�E�FPOS1 1�>��  x���� �Ώ���{���� :�Տ7�p����/��� S�ܟ���՟6�!� Z���~����=���د s����� ���D�V�� �=�����¿]�濁� 
ϥ��@�ۿd����� #ϬϾ�Y�kϥ���� *���N���r��oߨ� C���g��ߋ��&��� ���n�Y��-��Q� ��u������4���X� ��|���)�;�u����� ������B��?x �7�[��� ��>)b��! �E��{/�(/ �L/^/�/E/�/�/ �/e/�/�/?�/?H? �/l??�?+?�?�?a? s?�?O�?2O�?VO�? zOOwO�OKO�OoO�O �O_._�O�O_v_a_ �_5_�_Y_�_}_�_o �_<o�_`o�_�o�o|�2 1ш�2oDo~o �o�o &oD�oh e�9�]��
� ����d�O���#� ��G�Џk�͏���*� ŏN��r���1�k� ̟��🋟���8�ӟ 5�n�	���-���Q�گ u�����ӯ4��X�� |����;���ֿq��� ��Ϲ�B�ݿ��;� �χ���[����ߣ� �>���b��φ�!ߪ� E�W�iߣ����(��� L���p��m��A��� e����������� l�W���+���O���s� ����2��V��z '9s���� �@�=v� 5�Y�}��� </'/`/��//�/C/ �/�/y/?�/&?�/J? �/�/	?C?�?�?�?c? �?�?O�?OFO�?jO�O�O)O�O�o�d3 1ҵo_OqO�O)__ M_SOq__�_0_�_�_ f_�_�_o�_7o�_�_ �_0o�o|o�oPo�oto �o�o�o3�oW�o{ �:L^��� ��A��e� �b��� 6���Z��~������ Ə �a�L��� ���D� ͟h�ʟ���'�K� �o�
��.�h�ɯ�� �����5�Я2�k� ���*���N�׿r��� ��п1��U��y�� ��8Ϛ���n��ϒ�� ��?�������8ߙ߄� ��X���|����;� ��_��߃���B�T� f�����%���I��� m��j���>���b��� ��������iT �(�L�p� �/�S�w$ 6p����/� =/�:/s//�/2/�/�V/�/�O�D4 1� �O�/�/�/V?A?z?�/ �?9?�?]?�?�?�?O �?@O�?dO�?O#O]O �O�O�O}O_�O*_�O '_`_�O�__�_C_�_ g_y_�_�_&ooJo�_ no	o�o-o�o�oco�o �o�o4�o�o�o- �y�M�q�� �0��T��x���� 7�I�[��������� >�ُb���_���3��� W���{������ß�� ^�I������A�ʯe� ǯ ���$���H��l� ��+�e�ƿ��꿅� ϩ�2�Ϳ/�h�ό� 'ϰ�K���oρϓ��� .��R���v�ߚ�5� ����k��ߏ���<� ������5����U� ��y������8���\� ������?�Q�c��� ����"��F��j g�;�_��<�/45 1�?� ��n���f ���%/�I/�m/ /�/,/>/P/�/�/�/ ?�/3?�/W?�/T?�? (?�?L?�?p?�?�?�? �?�?SO>OwOO�O6O �OZO�O�O�O_�O=_ �Oa_�O_ _Z_�_�_ �_z_o�_'o�_$o]o �_�oo�o@o�odovo �o�o#G�ok �*��`��� �1����*���v� ��J�ӏn������-� ȏQ��u����4�F� X����ޟ���;�֟ _���\���0���T�ݯ x����������[�F� ����>�ǿb�Ŀ�� ��!ϼ�E��i��� (�b��Ϯ��ς�ߦ� /���,�e� ߉�$߭� H���l�~ߐ���+�� O���s���2���� h�������9�16 1�<����2� �������������� R��v�5� Yk}�<� `����U� y/�&/���/ �/k/�/?/�/c/�/�/ �/"?�/F?�/j??�? )?;?M?�?�?�?O�? 0O�?TO�?QO�O%O�O IO�OmO�O�O�O�O�O P_;_t__�_3_�_W_ �_�_�_o�_:o�_^o �_ooWo�o�o�owo  �o$�o!Z�o~ �=�as��  ��D��h����'� ��]�揁�
���.� ɏۏ�'���s���G� Пk������*�şN� �r����1�C�U��� �ۯ���8�ӯ\��� Y���-���Q�ڿu��� ��������X�C�|�� ��;���_����ϕ�����B���f�L�^�7 1�i��%�_����� ��%���I���F�� ��>���b����� ����E�0�i����(� ��L���������/ ��S�� L�� �l���O �s�2�Vh z�/ /9/�]/� �//~/�/R/�/v/�/ �/#?�/�/�/?}?h? �?<?�?`?�?�?�?O �?CO�?gOO�O&O8O JO�O�O�O	_�O-_�O Q_�ON_�_"_�_F_�_ j_�_�_�_�_�_Mo8o qoo�o0o�oTo�o�o �o�o7�o[�o T���t�� !���W��{���� :�Ï^�p������� A�܏e� ���$����� Z��~����+�Ɵ؟ �$���p���D�ͯh� 񯌯�'�¯K��o��
���yߋ�8 1� ��@�R���
���.�4� R��v��sϬ�G��� k��Ϗ�߳������ r�]ߖ�1ߺ�U���y� ����8���\��߀� �-�?�y�������� "���F���C�|���� ;���_����������� B-f�%�I ���,�P ��I���i ��/�/L/�p/ /�///�/S/e/w/�/ ?�/6?�/Z?�/~?? {?�?O?�?s?�?�? O �?�?�?OzOeO�O9O �O]O�O�O�O_�O@_ �Od_�O�_#_5_G_�_ �_�_o�_*o�_No�_ Ko�oo�oCo�ogo�o �o�o�o�oJ5n	 �-�Q���� �4��X����Q� ����֏q�������� �T��x����7��������MASK 1�û�����?XNO  ��~�MOTE  3�����i�_CFG ��p�����PL_RANGl�g�t��POWER ��õݠ|�SM_D�RYPRG %�p�%m���TAR�T �ծ#�UME_PRO������_EXEC_E_NB  d�x��GSPDX��������TDB��ϺR�M޿ϸI_AIR7PUR�� p�B�\<�ٛMT_�TР�n��OBOT__ISOLC1��8�蠥��9�z�NAM/E p�n�ۙ�OB_ORD_N_UM ?ը5��H844 �g��bҘ� ���/�(/�^/Ҧ�/���PC_T�IMEOUT�� �x�S232��1��4�γ L�TEACH PENDANPЅ��������l�j�M�aintenance Consg���߾�"��f�No Use���߮߀��0�B�T��h�N�PO2�RҤ�zz�e�CH_L[�3�p���	���?!UD1:���=R�VAIL��R�����x�e�PAC�E1 2�p�
 �濫��{鋓��⤢��9˺�8�?�%���%��� 4IDu������� Y������): !4�8�Uu��� ���/�):/ !/O/q���U/� ��/ ?�/?6??K? m//�/�/�/c?�/�/ �/�?O2O	OOi?{? �?�?�?_O�?�?�OGO _._@_'_eOwO�O�O �O[_�O�O�_o�_+_ <o#oQos_�_�_�_Wo �_�_�o�o8 Moo�o�o�o�o�o�o �D��4��I�k }���a���돀���0�B��+�X�2a�s�������W�͏ �����4�U�<�j�o�3~�������Ɵt� ���<���Q�r�Y���o�4������ѯ� ���)�8�Y��nϏ�vϤ�o�5��ʿܿ�  Ϯ�$�F�U�v�9ߋ��ߓ���o�6������ ����A�c�r��V� �������o�7��� �(�:���^�����@s���������o�8� !�3�E�W�{���������o�Gw �/ �m�
u d  /������ /Nl -S-L/�/p�d� z��/�/ �/�/??&?/./@. 1:n?�;�?�/�/(?�? �?OO*O<O2?D?V? h?�?�O�O�?�?HO_ _&_8_J_\_ROdOvO��O�O�_ ` @p��U]/o�O�IAakU�_Rodoj_Dj Eowo�o�o�o�o�o %�o�o=AS e���	���3� E���+�]���a�o\�
#o�o�_MOD�E  /
�S ��/㏙_�Z �oH�����	������CWORK_A�D�
����R  /< 1����_INTVAL��a�%�R_OPoTIONR� %����V_DATA_GRP 2�uX:D�@PП��̟ �˩͏���1��U� C�y�g�������ӿ�� ����	�?�-�O�u� cϙχϽϫ������� ���;�)�_�M߃�q� �ߕ߷��������%� �I�7�Y�[�m��� �����������E� 3�i�W���{������� ������/SA�we����P��$SAF_DO_PULS�Q�A���� CAN_TI�M��E}�R �� � �Ƙqsy�֡A��Yo�K�C կ ������l/�/%/7/I/[/e���C�2�$KKd��(�!�!ѢIf) �P5��/�/�/���)�/� ��4�_ �R  T0�!?^?�p?�?�9T D���?�?�?�?�? OO $O6OHOZOlO~O�O�O��O�O�OU�s��'��O$_6_�I  }�T;�o���WQo�p�M
�t��Di��[=Z0 � ��o�[Q [SC�_�_�_�_o  o2oDoVohozo�o�o �o�o�o�o�o
. @Rdv���� �����*�<�N� `�r��������?�� я�����+�=�O� ��r%{�������ß՟������"�_���0 2�SwU�]n������� ��ȯگ����"�4� F�X�j�|�������Ŀ ֿ�����0�B�T� f�xϊϜϮ������� ����,�>ߩ�b�t� �ߘߪ߼�������� o�(�:�L�^�p��� ���#�Q�[����
� �.�@�R�d�v����� ����������' 9K]o���� ����#5G Yk}�������O�3�//1/ C/U/g/y/�/�/�/�/��/�/�/	??-?;:p�D?q?{6��d��j?@]	123�45678�Rh!B!����B��V��?�? OO)O;OMO_OqOwA ��O�O�O�O�O�O_ _*_<_N_`_r_�_�_ �_�_�]�O�_ oo$o 6oHoZolo~o�o�o�o �o�o�o�o�_�_D Vhz����� ��
��.�@�R�d� #��������Џ�� ��*�<�N�`�r��� ������y�ޟ��� &�8�J�\�n������� ��ȯگ����ϟ4� F�X�j�|�������Ŀ ֿ�����0�B�T� f�%��ϜϮ������� ����,�>�P�b�t� �ߘߪ߼�{������ �(�:�L�^�p��� ��������� ����0.�@�%���l�~�����Cz  B}\�   ��}2d4� ���d1
���  	�d22,�%7I�Xp���Z�� ����� %7I[m�� ������!/3/ E/W/i/{/�/�/�/�/ �/�/�/??/?A?S?e?w?�?�:Z������<�4��`�$SC�R_GRP 1�� �  �� ߐ ��� ���	 �1��2
BD [����� I�7GDO2O�kO�����hBD?E� DP�wC��GhK�ARC� Mate 12�0iC 6789�0��M-�@A }8��M2IA�A���
12345t�D;F�2  ����>U�1{F�1HC�1��AhAJ<ANY	�?R�_�_�_�_�_�\��H��0�T�7�2 o/O0oVoho7F/��Co�o?o�o����l0Q�o:DBǲ�Ɛr2tAA��A c @��YuA@�WpNj ?�wrH����DzAF@ F�`�r��o��� ��B�-�f�Q���}�Yq�r������ďքB��y�*��N�9�r� ]�o�����̟���۟ �&���CTOF�k������h�����qYq6'���7G@Ypݯ����W\HC+�3���AnpC�V��o�~ec��W���  y���������ո�\�¿ P�(�@%�7�I�v�b�SS��0�EL_DEFAU�LT  m�����u�HO�TSTR��d���M�IPOWERFL�  ������W�FDO�� �� �u�RVENT 1����`�� �L!DUM_E�IPL�(��j!?AF_INE��Fߞ��!FT�u��<ߙ�!o�� ������!RPC_OMAIN���غ�ߜ1���VIS��ٻ� �}�!TPp�P�Ut�/�dl���!
�PMON_PROXY��2�e��������+�f�a�!R?DM_SRVb�/�9gP���!RT���0�h����!
��M�,�,�i��E!R�LSYNCFl	�84�!ROS�߸�4��!
�CE��MTCOMd�2�k�)!	�OCONS*1�l�u!�WASR�C|�2�md�!N�USB�0�n�>/!STM��'/.�o�Y/��}/p�J/�\/�/�/�/�/��ICE_KL ?%�� (%SVC�PRG1�/::$52�:???)03b?g?)04��?�?)05�?�?)06�?�?)07OO)0
T$JOE<9ROWK&4�� O)1,?�O)1T?�O)1 |?�O)1�?_)1�?G_ )1�?o_)1O�_)1DO �_)1lO�_Q1�OoQ1 �O7oQ1�O_oQ1_�o Q15_�oQ1]_�oQ1�_ �oQ1�_'Q1�_OQ1 �_wy1%o�/	2)0? "0��I1�/��S� >�w�b�������я�� ������=�(�a�L� s���������ߟʟ� �'�9�$�]�H���l� ����ɯ��ۯ���#� �G�2�k�V������� ſ���Կ���1���C�g�Rϋ��*_DE�V ���MC:��,�~��GRP 2�����0bx 	_� 
 ,���� ߟ���7��[�B�T� ��xߵߜ�������� ��3�E�,�i�P��� ����z��������� A�S�:�w�^������� ��������+O ��D�<���� ��'9 ]D ��z����� /h5/G/./k/R/�/ v/�/�/�/�/�/?? ?C?*?g?y?`?�?�? �?�?*/�?�?O-OO QO8OuO�OnO�O�O�O �O�O_�O)__M___ F_�_�?x_�_p_�_�_ oo�_7oo[omoTo �oxo�o�o�o�o�o �oE�_i{b� �������� A�S�:�w�^������� я�����^+��O� a�H���l�������ߟ Ɵ����9� �]�D� ����z�������� ���5�G�.�k�R��� ����ſ���������C�*�<�yϟ�d ���	gϰϛ��Ͽ�0�����+�%�+�P������i��i� y߇�qߧߕ��߹��� ��=�"�e���O�=�s� a���������3� ��'��K�9�o�]�� �������������# G5k�����[ �W���C �j�3���� ���/]B/�/ u/c/�/�/�/�/�/�/ 5/?Y/�/M?;?q?_? �?�?�?�/�?�?�?�? �?OIO7OmO[O�O�? �O�?�O�O�O�O�O_ E_3_i_�O�_�OY_�_ �_�_�_�_�_oAo�_ ho�_1o�o�o�o�o�o �o�oIooo@os a�����!� E�9��I�o�]��� �����ޏ������ 5�#�E�k�Y���я�� ����ן���1�� A�g�����͟W����� �ӯ	���-�o�T�f� �?���������Ͽ �G�,�k���_�M�o� qσϹϧ�����C� ��7�%�[�I�k�m�� ������ߥ����3� !�W�E�g���ߴ��� ���������/��S� ��z���C���?����� ����+m�R�� �s����� E*i�]K�o ����/A� 5/#/Y/G/}/k/�/� �/�/�/�/�/�/1?? U?C?y?�/�?�/i?�? �?�?�?�?-OOQO�? xO�?AO�O�O�O�O�O �O�O)_kOP_�O_�_ q_�_�_�_�_�_1_W_ (og_o[oIoomo�o �o�o	o�o-o�o!�o 1WE{i��o� �����-�S� A�w�����g�я�� �����)�O���v� ��?�����͟���ߟ �W�<�N��'��o� ����ɯ���/��S� ݯG�5�W�Y�k����� ſ��+�����C� 1�S�U�gϝ�߿��� �������	�?�-�O� ���Ϝ���u��߽��� ����;�}�b��+� ��'���������� U�:�y��m�[���� ��������-�Q��� E3iW�{�� �)�A/ eS����y� u�//=/+/a/� �/�Q/�/�/�/�/�/ ??9?{/`?�/)?�? �?�?�?�?�?�?OS? 8Ow?OkOYO�O}O�O �O�OO?O_OO�OC_ 1_g_U_�_y_�_�O�_ _�_	o�_o?o-oco Qo�o�_�o�_wo�o�o �o;)_�o� �oO������ �7�y^��'���� ����ُǏ��?�$�6� ���W���{����� ՟���;�ş/��?� A�S���w����ԯ� �����+��;�=�O� ��ǯ���u�߿Ϳ� �'��7ύ�����ÿ ]Ϸϥ���������#� e�J߉��}�ߍ߳� ��������=�"�a��� U�C�y�g������ ���9���-��Q�?� u�c������������ ��)M;q�� ��a�]�� %I�p�9� ������!/c H/�/{/i/�/�/�/ �/�/�/;/ ?_/�/S? A?w?e?�?�?�??'? �?7?�?+OOOO=OsO aO�O�?�O�?�O�O�O _'__K_9_o_�O�_ �O__�_�_�_�_�_#o oGo�_no�_7o�o�o �o�o�o�o�oaoF �oyg���� �'�����?� u�c���������#� ����'�)�;�q�_� ��׏�������ݟ� �#�%�7�m�����ӟ ]�ǯ���ٯ���� u���l���E�����ÿ ���տ�M�2�q��� e���uϛωϿϭ��� %�
�I���=�+�a�O� qߗ߅߻�����!߫� ��9�'�]�K�m�� �ߺ��߃�������� 5�#�Y������I�k� E���������1s� X��!�y��� ��	K0o�c Q�u����# /G�;/)/_/M/�/ q/�/�/�//�/? ?7?%?[?I??�/�? �/o?�?k?�?O�?3O !OWO�?~O�?GO�O�O �O�O�O_�O/_qOV_ �O_�_w_�_�_�_�_ �_oI_.om_�_aoOo �oso�o�o�oo�o �o�o�o']K�o ��o����� �#�Y�G�}����� m�׏ŏ������ U���|���E�����ӟ ������]���T��� -���u�����ϯ��� 5��Y��M�߯]��� q�����˿��1��� %��I�7�Y��mϣ� ���	ϓ�����!�� E�3�U�{߽Ϣ���k� ����������A�� h�z�1�S�-����������[�@�����$SERV_MA_IL  �����e�OUTPUT�t���RV �2�	�  �� �(�O���i�SAV�E��g�TOP10� 2�� d ��;M_q�� �����% 7I[m��� ����/!/3/E/ W/i/{/�/�/�/�/�/��/�/??/?	�Y�P��f�FZN_C�FG �	����.��o1GR�P 2�y7�� ?,B   A�0.�D;� B�0��  B4.R�B21��HELL�r2�	���������7"O1K%RSR 1O2ODO}OhO�O�O�O �O�O�O�O_
_C_._�g_R_�_�_�^�  ��%�_�_�_(�R�\a. �_b�`ރ��R2. d�o�_�6HK 1��; o�o�o�o �o�o�o�o
3.@ R{v��������<OMM ���?2��2FTOV_�ENBt����HO�W_REG_UI�R�g�IMIOFW�DL��!��5A���*SYSTEM�*. V8.303�40 ł11/9�/2020 Q� ���X�SN�PX_ASG_T�   0 $�ADDRESS � ��ZE�V�AR_NAM	��%$MULTIP�LY��PAR�AM�� � �$TIME����$�_ID�	$�NUM�D�T�CI{MP[�FRIFD�VERSION���G�TATU �$wDISK�NFOD��MODBUS_A�DR[�����POR�C���SSR~�� x ���NGLE��g�$�DUMMY7�S�GL�TASK   &����T�x�����STMTT0��PSEGT2�B�WD�h��E��SVCNT_GP��� 8 $PC��ER_V�  � 	$FB�PNm�SPC��m� S��DX�R[��� �$DATA0�Ӏ u���1��2���3��4��5��6���7��8��9��A*��B��C��D��2�B��F�� y���1ΩU1۩1�1��1�U1�1�1)�16�U1C�1P�1]�1j��1w�ҁJ���2Ω2�۩2�2��2�2��2�2)�26�2�C�2P�2]�2j�2�w�3��3��3Ω3�۩3�3��3�3��3�3)�36�3�C�3P�3]�3j�3�w�4��4��4Ω4�۩4�4��4�4��4�4)�46�4�C�4P�4]�4j�4�w�5��5��5Ω5�۩5�5��5�5��5�5)�56�5�C�5P�5]�5j�5�w�6��6��6Ω6�۩6�6��6�6��6�6)�66�6�C�6P�6]�6j�6�w�7��7��7Ω7�۩7�7��7�7��7�7)�76�7�C�7P�7]�7j�7�w�` ��PRM_�UPDӑ  s$4q� 
�����ӑؐ$TO�RQUE_CMDo   u�MOa�_SPEEjQ_�CURREo�nA�XI �mS�C�ART��_Uht��|P���LO�? � ��� ���������_�{�oVALU�OP���$�#(F�ID_�L��K%HIF*IN��$FILE_A�v$�$M�t���SAR0  h�^� E_BLCK����"���(D_CPU�)��)��F#y/�$����_=�R 	� � PWҐO�T��)1LA#�S�R� .3?184RUN_FLGQ5-4U184WITX5v1-4v185�H2�D4�084�TB�C2��
 � $O�X0IGu �0�_FTM1D��42�D�TDCX0AZ���2M���6�1�7THD��C�DxGR.0<A��ERVE�3?D��3?D3O��0_AC�@ X -$jALEN�3wD�3�j@EL_RATI6��$�W_�F#i1jAc$2�GMO�!�>��C��ERTIA��o!�Iaj@�KDE|�E��LACEM��CC�CmV�@MA���F7UW7QTCV8>\_QWTRQ^\U�uZ���Ct��USt�JI_��q�M�TF�J2'����E�QUvA2��P>�s�a�C@JKfVK�1'a�1'a`Af`J0<d+cJJ3c;JJ;cAAL+ca`(3ca`[f4\e5C�P�N1�\�`Q[;P�L��@_�E�W�3CF�� `^GRO�U1 ����y�N�0C�C��`REQUIR*B��EBUZ�fA�V7$T�@2#qg@pv�14 \��ENABL	�$oAPPRpCL��
$OPEN`xC/LOSEozSE�yr�E
�1.� �u �M�0<PPB�t_M	Gr!�pC��� �x���9P�wBRK�yNO�LD�vh�RTMO!_�3���uJ"��PcdP3cP;cPcP�cP6P��S�b���!�2�5� �r�B�1���1��PATH��ӁɃӁ�H�σ0�(p�W�SCaATr�ar�qINiB�UC�@��)�C��U%M2�Y�@+@�P9��O!EAT��0T�`@T�P�AYLOA�J2=L7R_AN�1���L*0���������uR_F2LSHR9DؑLO��(�ٗF��>F�ACRL_�!&���"���4bH$ ��$H�rG�FLEX�cs�1J�6 P@Mr�?�?>OPO� c�>iE :vO�F P٧�O5aP�O�O�LF1�>�R��O�O �O�O_!_��E+_=_ O_a_s_�_�_�_�_Y� vĽW�Sdf����_�_H o�jT2'W�X� `�eŴ��e'� �*o <oNo``deme[ee�oКo�o�i�2J�d ���0�o�o� 8A1Tk�q�PELٰ}1�=�xJ(p#pJE� �CTR"�f�TN�R9�wHAND_�VB�c�0 ��� $��F2�v	D6#SW�!�á�v� $$M�� �yv�q���q�����>��AR ���vQ!5���}A�| �zA�{A��@��{� �zD�{D��P�G@0��ST��w���y��N�DY W0^p�v!�H���k@ϗ �ϗꑎ�g������PX�a�j�s�|���p�����ӵ5 ���Ť����qAS�YM��^�p������_�0�.� A�+�-��K�]�o�����J��K�����˙.x�_VI��	(�s> V_UNIC.$P�בJeG"uG"� K$�X$|&
��P�K�,�>��%�T�\���2�0H+0Rr���!Lv�VrDI�sO4q�1� �c `�
O�I2AO�F�I1l��WW3o��1�۱�  � � ��M�E��@r2�"YT0PT���ڀ�1�`��du���8�1�9T���a $DU�MMY1`A$P�S_i�RF+�  tڀ�6XpFLA�`�YP��B�3$GLB_T��5*E�0�Vq�`��j�v1 XXMpw��ST±#p�SBR��M21_�VrT$SV_E�R��O� pC�CCL�D@pBAڰOL2� G�L EW� 4\�`�1$YQ�ZQ�!W�C`ԑ��As02�t-2�AU�E ��yN�@�$GIz�7}$�A �@�C�@� L�`V��}$F�EVNE+AR��Np�F]Y���TANCp��0�JsOG�A� ��$JOINT
Ѽ�`�EMSET��  WECU۱�S���!+Q���k g�U��?�#pLOCK_FO鐼��0BGLVm�G�LhTEST_X9Mcp�QEMP�Prq+bBB�P$U����B2�2#p�CQa�b���PQarACE��`Sr` $KAR��M3TPDRA8�@�d�QVEC��f֊PIUQaVaHE��PTOOL2��cVv1�RE�`IS3��r�b6s�f�ACH�P�(p�aO��3�42�9�2�`ISr  �@$RAIL_B�OXE
��@RO�BO"d?��AHOWWARO�Aq�0qROLM�2gu��
t�xr��/pZ���O_F��! ���@�a�] �_ �R�`Oˢ!!�r*��Q�p�Q�BKOU�R"XBMeY�C���P$PIP#fN���b/r�ax�Qa��p��CORDED��P��q� ��OY0 �# D )@OBu�G��Pd�S��3(@�S��I�SYSS�A�DRH�� �0TCHl�S� ,0EN2*�A�Q_T���Ѿ��PVWVAu1% � �`�B5PREV_RT��$EDIT�V/SHWR��\F$�����A	 D�0���;���$HEADД� U���KE|�A�0CPSPDl��JMPp�L5�3TR��44&[�t����I,`SH�C��N�E�`I��TICK�2�<M}����HNRA' @]����Վt�_GP�&v��S�TY��qLODA�P����m�( t 5
 �Gƅ%$�Tu=\@S>�!$=! 2��1EF0FP��SQU�`%�B!T�ERC�0��TS��) Ph@�� ����g��a�`O�0�3Ft�IZDQE�1�PRE��1!����pP9U�1�_DObR���XS�PK6AXI4P��sVaUR�ڳ@I�Hp�~����_�`��ET��P bl�%O�FP�AC�4 ss`�-2{SR��*lѠ ��A�������� #��1��A�R�c�R� s�RŃ�d�~Ͱ�dŢ� �����ː�C��|�����SC,@ o+ h�@DS�̐a�0SPC0~�AT�q��2�𐿒�2A_DDRES�cB��SHIF�H`_2+CHH�z�IK@��W�TV�I72,��Ph���� 
+j
�rqV�qA���- \�����O����<�C���򢵲���B<��TXSCREEU��.	0k�TINA�CP��T�Q����� / T���@��� �Ag@��^���^����RROL wP��f����v�-1UE��0 ��� ��@S�A��RSyM�T�UNEX��6F�� S_�Cf�6 V�i���6��C�RB���� 2/��UE��1=2�B��!�GM�T� Li!m�w@O^�WBBL_pW�0N��2 �O�O�A�LE��GpTyO�3RIGH&�BRD�D��CKG9R�0NTEX��O>JWIDTHs1��u�"qA�a%�I_��0H�� 3 8��!wP_T��ҭ�0R��@�Rsw�2$� O��ѭ�4���GG U�2 �R brqLUM8�u���ERV
��@�� PaP�У5{0^�GEUR&cF����Q)]�LPM��E��C�)jS�x�xT�`w5u6u7u8Z���3�9P��6j�a�QS��4��USR�D6 <ĥ��0UR��RFO�C�aPPRIαmxp�!L TRIP+q�m�UN$0547	Pt�$0��Yq5%�8Ia���� 8� . �G \�T�p1�L�ѣ"OS�1�&R���#�a�9�O�C�N��"�$�IaUU�:��/�/�U��#OF�F!`��;[�3O�n0 ٰW5�4:N�@GUNw��0B_SUB�2p@��'SRT� �<��vQ̗p �ORp�5RA�U��4T�9���1_����= |���O�WN� T$SRC���r�D!`CEMPFI*�*ё�ESP-������e*B��&�b�!B���> M`10WO8�T�n��COP:1$���� _^@�b�A�q�EWA�C?a�A�@�C�A>�C �VCCH��? �qC36MFB1�%R4�Y`��@x %rT���AXdP^��spC�p^RUDRIV���C_V�uT̐fpD�?MY_UBY�ZT V�񕠧�B��X�a��RP_Sp�+��RL�7�BM$��DEY��EX����E�MU��X7d[�UASP�po��G���PACINΑ}�RGMAadwbF3wb3wb���ARE����a�r#7Swb�pA R�@EG�PPr�`5VR� �pB d�_���2�	�BN�RECcSW&o`_Apa�8c��O!��A��1s�E��UB�� �q5VHKG�C��Iz���.p��zsEA���w�@x� 1u5UMRCV��WD �FOS�M� �Cs�	�rX3�c�rREF���v�v�q p7 ��p �z��z��{;��vp_@@�zq��{��S�/g�Sᡏ�#�8R��E �$�=�hߠ) �UӠOU�x�b�ZS @�e
2�2�$��R� �ΐ�B��2Ѻ�Kq�S�ULs�C�@CO�:�� D)`�NT �CZ��BY��e�!e�$�L�S���S������!�JTǤFt� +��ǱT� ��C7ACH+�LO�����*`����@ܣC_oLIMI��FR%�qTj�'���$HO� z6B�COMMpSB�O0 ]�Ԉ�I؄�h@VP�b��_S�Z3n���6����12���[`��&����AvaMP�FAI&�5Gvt��AD��B�MREׄ9�_SI�Z�PH�`��FA�SYNBUF�FV�RTDk�w�I�aOML��D_@3��W3�P�ETUc�Q�Np[�ECCU�hV�EM�`��۲&�VIsRC���VTP�p�O��J�s�A�w�_DGELA�cP�ƫ�`�KS��G�@9pCKWLAS�3	ő_�$F�ƀHp"�S;��yN��PLEXEE�I��B/��3cFLK I `]�^A��M���dws��/�^@�bJ# �ʱ��#�#\RS ORD@!�4QP> 3 ނ)�K���T\"���WwCb2V��g%L`�Qۑ6D�4��\*bUR3cp_R'�d���,a]��ծc �_od&�{g��`Br*�T�'�SCO��*�C� ad�"_f�"0� �">�"K�"Y�J_\_�nZ��� E\ AMܐP�0 PSM�f%Mp"%HADJ�T�/e��Bڒ� N8p"q׬!LIN]3q�/�XVRh$O\����T_OVR� �/ZABC�5P�bw�t$��
4QZIPg%}Qp"DBGLV�C�L�R ��J�ZMwPCF�5R  r ����$��QLNKʦ2
u�M,a|�S ��|q����CMCM�i`C�CC�ACtP�_�  $J:4D��@QJ��V�4$0�tO�UsXW� ��UXE>a ��E�[���	��u��T P����r�YK�D"0� U�"��^I3GHbcq�?( �K���V � vG��$B$��@1e��B�҉�&GRV%�F8� ���OVC�5@�A7�w@�`��
VB�I���D�TRA�CEB�V�1�SP�HER�P W �, �3I[�$S�IM�A�!2Re!� ��e!V&��qe!q�m/!��%���/8Kpb/t#_UN�@_+7p&LCд�%� �%V M��A�LIAS ?e����%1�! ( he�!:?L?^?p? �?�66?�?�?�?�?�? 	OO-O?OQO�?uO�O �O�O�OhO�O�O__ )_�OM___q_�_._�_ �_�_�_�_�_o%o7o Io[ooo�o�o�o�o ro�o�o!3�oW i{�8���� ���/�A�S�e�� ��������я|���� �+�֏<�a�s����� B���͟ߟ����'� 9�K�]�o�������� ɯۯ�����#�5�� Y�k�}�����L�ſ׿ ���ϸ�1�C�U�g� y�$ϝϯ�����~��� 	��-�?���c�u߇� �߫�V��������� ��;�M�_�q��.�� ���������%�7� I���m��������`� ������!��EW i{&����� �/AS�w ����j��/ /+/�O/a/s/�/0/ �/�/�/�/�/�/?'?�9?K?]?3�$SM�ON_DEFPR�O �����1 �*SYSTEM*�p:RECALL �?}�9 ( �}d?�?�?�?OO0O �?UOgOyO�O�O�O BO�O�O�O	__-_�O Q_c_u_�_�_�_>_�_ �_�_oo)o�_Mo_o qo�o�o�o:o�o�o�o %�oI[m ��6������!��~*copy �mc:diocf�gsv.io m�d:=>172.�8.9.225:142242���������z4F�frs:�orderfil�.dat vir�t:\temp\@]�o�
��.��q,Ɔ*.dڏ�󏄟������w
xyzra?te 11 Q�c� u���*��uƗߟ4 ����������t�7Ə؈mpbac�kޟx���0� }-.F�dbN�*ۯ�`���������u2xƤc:\O�аa�4 y�P
��.��q3Ƶaο �n����Ϟϰ�ïկ ^���
��.�A���e� �ψߚ߬߿�R�d��� ��*�=�����sτ� ������V����� &�9�K���o߀����� ����\�����"5� G���k�2��3ř�Qcu*�u<F���8644�� ������Qcu�//*/=�O�0836 ���/�/�/�� ��Y�Z'�/?!?4�F� �/Y(�/�?�?�?=�/<؏��680 z?OO/O� +F��?�5�? �O�O�O:L/mCdOvO�__+_�$:�4h:�\support�PPY=>4798�54592:64327�O�_�_5_G��TCoutput\�untitled�8.pcY� overm__o"o�_�_�T9�_�_�o�o�o�'�tpdisc 0�O aoso(��'tpconn 0��o�o2����{�$SNPX_�ASG 2 �����q�� P 0 '�%R[1]@1�.1��y?��#% �(��L�/�A���e� ������܏��я��� �H�+�l�O�a����� ��؟����ߟ�2�� <�h�K���o���¯�� ̯��ۯ����R�5� \���k��������ſ ����<��1�r�U� |Ϩϋ��ϯ������ �8��\�?�Qߒ�u� ���߫�������"�� ,�X�;�|�_�q��� ����������B�%� L�x�[���������� ����,!bE l�{����� �(L/A�e ������/� /H/+/l/O/a/�/�/ �/�/�/�/�/�/2?? <?h?K?�?o?�?�?�? �?�?�?O�?ORO5O \O�OkO�O�O�O�O�O �O_�O<__1_r_U_ |_�_�_�_�_�_o�_ o8oo\o?oQo�ouo�o�o�d�tPARAoM �u�q_ �	��jP;tUAp�h#t��p�OFT_KB_CFG  s�u�s�OPIN_SIM  �{vu���p�pRVQST_P_DSB^~r���x�`SR >ay � &(u��#��vTOP_O�N_ERR  �"uJy?�PTN z�fr�A;��RING_PRM�I� �`VCNT?_GP 2au&q�(px 	�̏p`���ޏ��wVD���RP 1�i'p �y�R�d�v����� ����П�����*� <�N�`����������� ̯ޯ���&�M�J� \�n���������ȿڿ ���"�4�F�X�j� |ώϠϲ��������� ��0�B�T�f�xߟ� �߮����������� ,�>�e�b�t���� ���������+�(�:� L�^�p����������� ���� $6HZ l~������ � 2DV}z �������
/ /C/@/R/d/v/�/�/ �/�/�/�/	???*? <?N?`?r?�?�?�?�?��?�?�?OO&O0�P�RG_COUNT�?v�r�NuRBEN�B��MEMwCAt�O_�UPD 1�{T  
;Or�O�O �O__(_:_c_^_p_ �_�_�_�_�_�_�_ o o;o6oHoZo�o~o�o �o�o�o�o�o  2[Vhz��� ����
�3�.�@� R�{�v�����Ï��Џ ����*�S�N�`� r����������ޟ� �+�&�8�J�s�n��� ������ȯگ���� "�K�F�X�j������� ��ۿֿ���#��0��B�k�f�x�DL_IN�FO 1�Es�@��	 ����������@L�g�@�D�?���{�	
� ��	̀��@������%^���A�f���o߁� D���D�q}D�Q�6��p´�����O@YSDEBU)G\@�@��d�I��SP_PASS\E�B?��LOG ����C����ؘ�  ��A��?UD1:\���_MPC�E��$��AH�� �Am�?SAV �m��4�L��S�SV�d�TEM_TIM�E 1	��@+ 0������_���$T1SVGU�NS�@]E'�E��r�ASK_OPT�ION\@�E�A�A���_DI��xO��B�C2_GRP 2�
�I=���Ѡ  �C�f�BCCF�G ���� l�]`]`ߕ ������� 7"[FX�|� �����/3// W/B/{/f/�/�/�/�/���,�/�/"?4?�/ ?j?U?�?y?�?���? ���0�? O�?$OOHO 6OlOZO|O~O�O�O�O �O�O_�O2_ _B_h_ V_�_z_�_�_�_�_�_ �_�_.oh� BoToro �o�oo�o�o�o�o�o &8\J�n �������"� �F�4�j�X�z����� ď���֏����� 0�f�T���@o����ҟ ���t���*�P�>� t�����f������ί ����(�^�L��� p�����ʿ��ڿ �� $��H�6�l�Z�|�~� ���ϴ��Ϡ���2� D�V���z�hߊ߰ߞ� ���������
�@�.� d�R�t�v������ �����*��:�`�N� ��r������������� ��&J �bt� ��4���� 4FX&|j�� �����//B/ 0/f/T/�/x/�/�/�/ �/�/?�/,??<?>? P?�?t?�?`�?�?�? OO�?:O(OJOpO^O �O�O�O�O�O�O _�O $__4_6_H_~_l_�_ �_�_�_�_�_�_ oo Do2ohoVo�ozo�o�o �o�o�o
�?"4R dv�o����� ����<�*�`�N� ��r�������ޏ̏� ��&��J�8�Z���n� ����ȟ���ڟ���� �F�4�j� ������ į֯T����
�0���T�>�r��$TBC�SG_GRP 2�>�� � �r� 
 ?�  ������ӿ ������-��Q�c��v�}���d0� ���?r�	 H�C�`�r���b�C�  B����Ȟ��>�ff�źƞH�������϶�\���H �h�BLcφ�B$дh�j߈ߎ߰�H�����ތ��@�@�� AƷ�f�y�D�V����������	��?33�3��2�	V3�.00��	m2;ia�	*T�L�pq�c�"����r����� ��l���_   ��B��X����u�J2}����5���CFG ->��� ��
��D��o�o��
G���� ���5 YD V�z����� �/1//U/@/y/d/ �/�/�/�/�/�/�/? ???Q?����\?n?�? *?�?�?�?�?�?O�? 1OOUOgOyO�OFO�O �O�O�O�O	_r�^�._ :�>_@_R_�_v_�_�_ �_�_�_�_o*ooNo <oro`o�o�o�o�o�o �o�o8&\J l�������� ���6�X�F�|�j� ����ď��ԏ���� ܏.�0�B�x�f����� ��ҟ�������*� ,�>�t�b��������� �ί���:�(�^� L���p�������ܿʿ  ��$��H�6�X�~� (��ϨϺ�d������� ���D�2�h�Vߌߞ� ���߀�����
���� @�R�d��t���� �����������*� `�N���r��������� ����&J8n \~������ "��:L
� |������� 0/B/T//d/�/x/�/ �/�/�/�/?�/,?? P?>?`?�?t?�?�?�? �?�?�?OOOLO:O pO^O�O�O�O�O�O�O �O_ _6_$_Z_H_j_ l_~_�_.�_�_�_�_  oo0oVoDozoho�o �o�o�o�o�o�o
 @.Pv��Tf ������<�*� L�r�`���������ޏ ̏����8�&�\�J� ��n�������ڟȟ�� �"��F�X�op��� o>�į���֯��� �B�0�f�x���H�Z� �����ҿ��,�>� ��b�P�r�tφϼϪ� �������(��8�^� L߂�pߦߔ��߸��� ����$��H�6�l�Z� ��~�������d��� �&�����D�V���z� ����������
. ��R@bdv�� ����*N <^`r���� ��//$/J/8/n/ \/�/�/�/�/�/�/�/ ?�/4?"?X?F?|?�? 8��?�?�?t?�?�?O O.O0OBOxOfO�O�O �O�O�O�O�O__>_�(^  dPhS �hV|_hR�$TB�JOP_GRP �20U��  ?�hV	��R�S�\�8P���p���Q�U  � �� � ��RhS �@dP�R	 �C�� ff  Cq�W�Q4b��<f>9o >�ff\a<a�=�ZC�`����b�&`H&`.g�o�gnѴW4e\e�`b�o ?a�d=�o7LC�noBȂo�#&`�`9u�o�c��33\uX2h�P<���C\vc@333@33|b}`f�BL�wHqDa�l����u�Jh�p�<X��B$�d���?���C*p��C���Z`y�<x��k< ��q`?]`C4.�ϏR�d��daG����{�<g���]p@&b`yap�c�z{ 4ep�V���������� ʟ���(�� �N�� Z����������ޯ�ʢd�hV0�4e	�V3.00�Sm72ia�T*Z��T�cQh�s� E��'E�i�F�V#F"wqF>���FZ� Fv��RF�~MF����F���F���=F���F��ъF��3F����F�{G�
GdG��G#
��D���E'
E�MKE���E��ɑE�ۘE���E���F���F��F���F(��F�5��FB��F�O��F\��F�i��Fv��F���vF�u�<#�
<t���	@Ť�r_X�j�M��hTn�@�U�S��SE?STPARSA�\X�P�SHR��ABL/E 1�[��hS��ȃ� �0cɞ�B����gWoQ��	��E
������hQ�������C���RD	I�ϬQ��� �2�D�Vվ�O�������ߐ��*���S�ߪS  �������!�3�E�W� i�{������������� ��/A�]���� �̂	k�}���M�_��q߃ߕߧ���hNUoM  0U�Q�PpP B�C���?_CFG P��a@�PIMEBF_TT����S���GVERAÔ���R 1�[ 8Ie�hRcP! 3P�  � //$/6/ H/Z/l/~/�/�/�/�/ �/�/�/? ?2?{?V? h?�?�?�?�?�?�?�>��?O�:0OBOTO .OxO�OdO�O�O�O�O �O�O_,__P_b_�8�_�_�_~_�_�_�_H�_���_K�@����MI_CHA�N� � mcDB'GLV逡����p`ETHERADW ?���`�n���?o�o�o��p`R�OUT�!p
!�"t@|SNMA�SK�h��a255.~uF�|��F����OOLOFS_�DI��GT �iO�RQCTRL Ip	��n��T� B�T�f�x��������� ҏ�����,�>�P��b�r����������PE_DETAI�h��zPGL_CON?FIG Qa���/cell�/$CID$/grp1��3�E�W�i�{�1�	����ʯܯ � ���$�6�H�Z�l� ~������ƿؿ��� ����2�D�V�h�zό� ϰ���������
ߙ� .�@�R�d�v߈��)߀����������} ��N�`�r��������턬���)� ;�M�_��߃������� ����l�%7I [m������� �z!3EWi �������� �///A/S/e/w// �/�/�/�/�/�/�/? +?=?O?a?s?�??�? �?�?�?�?O�?'O9O KO]OoO�OO�O�O�O��O�O�O_���User Vie�w !�}}1234567890B_ T_f_x_�_�_�T-`��_��(Y25Y�Oo o*o<oNo`o�_�_/R3�_�o�o�o�o�ogo)�^4�obt�@�����^5Q �(�:�L�^�p�����^6�ʏ܏� ��$���E��^7��~��������Ɵ؟7����^8 m�2�D�V�h�z��������� l?Camera3Z)�����(�:�L�*�E �v�����@_��ƿؿ0�����  ̦�Y �^�pςϔϦϸ�_� ���� �K�$�6�H�Z�l�~ߥ��̦�i��� ���� ��$���H�Z� l�ߐ��������� �ߣ�Py��6�H�Z�l� ~���7������#���  2DV���*� ���������� "4F�j|�� ��kͥ��Y/ / 2/D/V/h/�/�/�/ ��/�/�/
??.?� ��l��/z?�?�?�?�? �?{/�?
OOg?@ORO dOvO�O�OA?�� �1O �O�O
__._@_�?d_ v_�_�O�_�_�_�_�_o�O�G9�_GoYoko }o�o�oH_�o�o�o�_ �o1CUgy�	Υ0�o���� ���o2�D�V��oz� ������ԏ{�Ӡ իx�-�?�Q�c�u��� .�����ϟ���� )�;�M��ΥA�䟙� ����ϯ�󯚟�)� ;���_�q��������� `��u��P���)�;� M�_���ϕϧ���� ������%�̿޵� ��q߃ߕߧ߹���r� ����^�7�I�[�m� ��8�޵�(����� ��%�7���[�m�� ��������������� ޵���I[m� �J����6!�3EWi  	�������//(/:/L/^+   nv�/�/�/�/ �/�/ ??$?6?H?Z? l?~?�?�?�?�?�?�? �?O O2ODOVOhOzO �O�O�O�O�O�O�O
_ _._@_R_d_v_�_�_p�_�_�_b,  
 �(  �( 	 �_oo:o(o ^oLo�opo�o�o�o�o��o �o$�Z~* ̸i{� � �����X5� G�Y��}�������ŏ ׏�����f�C�U� g�y��������ӟ� ,�	��-�?�Q�c��� ������������ �)�;���_�q���ʯ ����˿ݿ��H�%� 7�Iϐ�m�ϑϣϵ� ��� ����!�h�E� W�i�{ߍߟ������� ��.���/�A�S�e� �߉����������� ��+�r��a�s��� �����������J� '9K��o��� ����X5 GYk}���� ��0//1/C/U/ g/��/�/�/��/�/ �/	??-?t/Q?c?u? �/�?�?�?�?�?�?:?p@ B"O4OFO�CG `��)f�rh:\tpgl�\robots\�m20ia\ar�c_mate_1>�@c.xmlO�O �O�O�O�O__(_:_L_XX��X_}_�_�_ �_�_�_�_�_oo1o CoZ_Toyo�o�o�o�o �o�o�o	-?Vo Pu������ ���)�;�RL�q� ��������ˏݏ�� �%�7�N�H�m���� ����ǟٟ����!� 3�J�D�i�{������� ïկ�����/�F� @�e�w���������ѿ������+�=�_HΕ1 Oj@88�?�=�|�=� xϚϜϮ�������� 0��<�f�P�rߜ߆�����߼����&��$�TPGL_OUT?PUT "H1H1_ `�H� ]�o��������� �����#�5�G�Y�k� }����������������H�`���2345?678901 2 DVhz�>2� �����9 K]o�}�� ������1/C/ U/g/y/�/#/�/�/�/ �/�/	?�/???Q?c? u?�??1?�?�?�?�? OO�?%OMO_OqO�O �O-O�O�O�O�O__ �O�OI_[_m__�_�_ ;_�_�_�_�_o!o�_ /oWoio{o�o�o7oIo �o�o�o/�o= ew���E��@���+�� �}[��a�s���������̍@�b����h� ( 	 7�%�[�I� �m���������ǟ�� �!��E�3�i�W�y� ����ï���կ������/�e�S���� ^�w���ѽ���� �)�;���d�v�� �Ϭϊ�����L���� ��(�N�,�>߄ߖ� � ����n������&�8� ��D�n��^���� ����V��"���F�X� 6�|�����z�����x� ����0B��fx �����N` ,�Pb@�� ��p�/�/ :/��p/�/$/�/�/ �/�/�/X/�/$?�/4? Z?8?J?�?�??�?�? z?�?O�?2ODO�?PO zOOjO�O�O�O�O�O bO_._�OR_d_B_�_ �__�_�_�_�_oo��_<oNoTb�$TP�OFF_LIM ����p�����qibN_SVm` � ӄjP_M�ON #����d�p�p2ӅiaS�TRTCHK �$��f^��bVT?COMPAT�hq��fVWVAR �%�mAx�d R�o Y�p�bia�_DEFPROG 3vb%p��d�_DISPLAY�t`�n�rINST_�MSK  �| ��zINUSER��tLCK��{QUICKMENA���tSCRE`����rtpsc@�t�{���b��_���STziRACE_CFG &�i�Atx`	bt
?��܈HNL 2'"�i}� �H{ nr4� F�X�j�|�������Ě�ޅITEM 2(� � �%$12�34567890<��  =<�7�<I�Q�  !W�_�kp���bs�ů)� ���_������^��� y�ݯ����5�%�7�I� c�m�翑�=�c�u�ٿ �����!ϛ�E���� )ߍ�5߱�����Yߧ� �����A���e�w�@� ��[�����ߧ�� k���O��s��E�W� ��c������}�'��� ��o�/������; S����#�GY "}=�as�� ��1�U/'/ ������_/	/ �/�/�/Q/?u/�/�/ ?�/i?�?�??�?)? ;?M?�?O�?COUO�? aO�?�?�OO�O7O�O 	_mO_�O�Ol_�O�_ �O�_�_�_3_�_W_i_ {_�_�_Koqo�o�_�o oo/o�o�oeo%7 �oC�o�o��o� ��O�s�N�ڄ�S�)�S�� 3 ϒS� �����y
 ��ݏď�~��UD1:\����e�R_GRP� 1*��� 	 @�pY�k�U�@��y�����ӟ���� ���͑�2��V�A�?�  q���m��� ��ǯ���ٯ����� E�3�i�W���{��������	!����c��SCB 2+o� \�Y�k�}Ϗϡ���������Y�V_C�ONFIG ,�o�󁧏�M���OUTPUT -o�>���Yߝ߯� ��������	��-�?� Q�c�u�;ъߝ���� ������	��-�?�Q� c�u������������ ��);M_q �������� %7I[m� ������/!/ 3/E/W/i/{/��/�/ �/�/�/�/??/?A? S?e?w?�/�?�?�?�? �?�?OO+O=OOOaO sO�O�?�O�O�O�O�O __'_9_K_]_o_�_ �O�_�_�_�_�_�_o #o5oGoYoko}o�_�o �o�o�o�o�o1 CUgy�'�9Ո� �����#�5�G� Y�k�}������oŏ׏ �����1�C�U�g� y���������ӟ��� 	��-�?�Q�c�u��� ������ϯ���� )�;�M�_�q������� ��˿ݿ���%�7� I�[�m�ϑϣϴ��� �������!�3�E�W� i�{ߍߟ߱������� ����/�A�S�e�w� ������������ �+�=�O�a�s����� ����������' 9K]o���� �����#5G�Yk}����x������� /�3/E/W/i/{/�/ �/�/�/�/�/�/?� /?A?S?e?w?�?�?�? �?�?�?�?OO*?=O OOaOsO�O�O�O�O�O �O�O__&O9_K_]_ o_�_�_�_�_�_�_�_ �_o"_5oGoYoko}o �o�o�o�o�o�o�o 0oCUgy�� �����	��, ?�Q�c�u��������� Ϗ����(�;�M� _�q���������˟ݟ ���%�6�I�[�m� �������ǯٯ��� �!�2�E�W�i�{��� ����ÿտ������,��$TX_SCREEN 1.����}�ipnl/`�g?en.htm,����ϣϵ���$ P�anel setup��}�����0�B�T�f����ϝ� ����������n��� ?�Q�c�u����"� ��������)����� ��q�����������B� ��f�%7I[m ���������� t��EWi{� ��:��//�//A/�/�UALR�M_MSG ?L��Y� Z//��/ �/�/�/�/�/??$? B?H?y?l?�?�?�?u%�SEV  �-��6s"ECFG �0L�V�  }/�@�  A#A�   B�/�
 �?6�L�VOhOzO�O �O�O�O�O�O�O
_W~�1GRP 21	Kw 0/�	 @O�b_u I_BBL_NOTE 2	J�T��l�6�Q�8�@uRDE�FPRO %�+ (%�?�_8��_o �_'ooKo6oooZo�o��o�o�o�o�ok\INUSER  �]�P_�oI_MENH�IST 13	I � ('p ���(/SOFTP�ART/GENL�INK?curr�ent=menu�page,153�,17������)q�~381,23�/�A�S��p�195���ԏ��p'y��4��3�E� W�i��q�o������ǟ ٟ�z��!�3�E�W� i���������ïկ� v����/�A�S�e�w� �TEplq�����Ϳ߿ ���'�9�K�]�o� ��ϥϷ��������� �Ϡ�5�G�Y�k�}ߏ� ߳����������� 1�C�U�g�y���,� ��������	����?� Q�c�u����������� ����),�M_ q���6��� %7�[m ���D���/ !/3/�W/i/{/�/�/ �/�/R/�/�/??/? A?�/e?w?�?�?�?�? �����?OO+O=OOO R?sO�O�O�O�O�O\O �O__'_9_K_]_�O �_�_�_�_�_�_j_�_ o#o5oGoYo�_}o�o �o�o�o�o�oxo 1CUg�o��� ����?�?�-�?� Q�c�u�x������Ϗ �󏂏��)�;�M�_� q��������˟ݟ� ���%�7�I�[�m�� � ���ǯٯ���� ��3�E�W�i�{�������ÿտ��������$UI_PAN�EDATA 15����A��  	�}�/frh/cgt�p/wholed?ev.stm�{���ϟϱ���)prii��ϧ�}���"�04�F�X�j� )lߐ� wߴߛ���������� 2�D�+�h�O�������� �    xh�����#�5�G� Y���}��ϡ������� ����b�1U< y�r������	�-?&c��  D��CÞ����� ��P!/��E/W/i/ {/�/�//�/�/�/�/ �/?/??S?:?w?^? �?�?�?�?�?�?Oz �=OOOaOsO�O�O�? �O./�O�O__'_9_ K_�Oo_V_�_z_�_�_ �_�_�_o#o
oGo.o ko}odo�oO&O�o�o �o1�oUg�O ������L	� �-�?�&�c�J����� ��������ڏ��� ;��o�o~�������� ˟ݟ0��t%�7�I� [�m��柣�����ٯ �������3��W�>� {���t�����տ�Z� l��/�A�S�e�w�ʿ ������������� +ߒ�O�6�s�Zߗߩ� ���ߴ������'�� K�]�D����Ϸ��� �������d�5�G��� k�}���������,��� ��C*gy `����������}�,ew����)S�W� �/"/4/F/X/j/� �/u/�/�/�/�/�/? �/0?B?)?f?M?�?�?��?�?Q�����$U�I_POSTYP�E  ��?� 	 �?#O��2QUICKME/N  KO&O��0RESTORE� 16��?  ��?X�!�O�C�OX�m�O�O __'_9_�O]_o_�_ �_�_H_�_�_�_�_o �Oo0oBo�_}o�o�o �o�oho�o�o1 C�ogy���Zo ���R�-�?�Q� c����������Ϗr� ���)�;����Z� l�ޏ����˟ݟ�� ��%�7�I�[�m���� ����ǯٯ�����
� |�E�W�i�{���0��� ÿտ���Ϯ�/�A��S�e�w�1GSCRE�A@?FMuw1sc�@u2��U3��4��5��6���7��8���2USE�R���ϫ�T����k�s���4�5�6��7�8��0ND�O_CFG 7�K<;�0PDAT�E ������ޝ4B��_I�NFO 18����RA0%}���Q��� �����'�
�K�]�@� ��d������������*L��OFFSE/T ;FM�� �@ �b�t��������� ������N�UL ^��������&VO(
L*�U�FRAME  ��d֑�RTOL_ABRTp�ӈ�ENB��GRP� 1<�IRACz  A����� �	//-/?&I/[/Ā@@U�iѠMS�K  ��ӢNm%��%��/�O_EVN��$c֬
6U�2=I9h�i�UEV�!�td:\eve�nt_user\��/T0C7Y?)�F��<L1SPR1W7spotweld�=!C6�?�?�?�@�$!�/h?&O[OGl� OJO8O�O�OnO�O�O �O_�O�O�Oe__�_ 4_F_|_�_�_�_�_�_ �_=o,oaooo�oBo �o�oxo�o�o'�o��j)6WRK 2>�@�88"��  y����
��.� @��d�v�Q������� Џ⏽����<�N��)�_������$VC�CMU�?\ݨ�MmR�2E8;<Ԝ"�	j���~?XC56 *�����h� �5�Vi�A@7 p? ȗ�' ;[�e�Ȁ����ů����^�9%A��ٯ*�� B���E� �I�ѯj�����]��� ��ֿ�������0χ� �f�Q�cϜ�O��������ISIONTM;OU? ��ů��FU��U��(� FR:�\��\u�A�?  �� MC*��LOG7�   7UD1*�EX[�E!�' B@ ����o�r���o�������d �  =�	 1- n?6  -������6,�ր�1�=�̩�:���n�P�TRAIN����1�E!��Ad��͓G8; (��:��S����� ������-��1�?�Q��c�u�������T���_��RE��H�����/LEXE��I8;��1-e��VMPH?ASE  ����A���RTD_F�ILTER 2J.8; ��R�� �����1 C#��t��������//��SH�IFT�"1K8=<a���/p/3��O/ u/�/�/�/�/�/�/? �/?)?b?9?K?�?o?��?�?�?	LIV�E/SNAP�3?vsfliv4�?���� SETyU�0BmenuO�O�?}O�OfB/%L���	|H{O�O�ô?�J� �@-�AVdB8�����K�HM�QR�S����	'-_ME�0�ļ��/!MOM ��zWqWAITDINEND����TOK  噰\��r�_S�_�YTIM����
lG�_,m�_�Ok�_/j�_/jo�XRELEK_g���Q��<֗Q_ACT�0^ht(q�X_3� N���)r%�O_��rRD�IS�0�n�$X�VR�BO �$Z�ABC͒1P��� ,����2g7Z+IP�CQ����/��A�S��zMPCF_OG 1R�J�0�X�w��a�MP�sS����<�����8�����3�̟�?�  �����̟ȿ������D���D�q}D��Q���?����:��hK=�&�7��);��=>�T�d��(�:�;B�T�f�v�e�Ο�����A�2�6��p´$�6�>Ȇ�n� h�z�����ȫ�pt���T|��w�YLIN5DqU|�  �e� ,(  *)��:���&�c�J���n� ���Ͽ�#��s� (��!�^ϡ��ϔϦ� ���e�K� ���$��`y�Z�l��{��2V�+q đ������ �������٧�D����^�A���SPH�ERE 2W	�� �Ϛ�ߓ������<� O�*�<���`������ }��������I�[� 8��\CU��������pZZ�f � �f