��   b�A��*SYST�EM*��V8.3�0340 11�/9/2020 A   ����CELLSE�T_T  � w$GI_ST�YSEL_P �7T  
7ISO:iRibDiTRA�R|��I_INI; �����bU9A�RTaRSRPNSS1Q23U4567y8Q
TROBQ?ACKSNO� �)�7�E� S�a�o�z�2 3 4 5* 6 7 8aw.n&GINm'D�&� �)%��)4%��)P%���)l%SN�{(O�U��!7� OPT�NA�73�73.:BP<;}a6.:C<;CK;�CaI_DECS�NA�3R�3�TR�Y1��4��4�PTHCN�8D�D>�INCYC@HG��KD�TASKOK�{D�{D�7:�E �U:�Ch6�E�J�6�C�6U�J�6O�;0U��:IATL0RHaRbH<aRBGSOLA�6�VbG�S�MAx��Vp��Tb@SEGq��T��T�@REQ �d�drG�:Mf�G�JO_HFAUL��Xd�dvgALE@� �g�c�g�cvgE� x�H�dvgNDBR�H<�dgRGAB�Xt�bT  �CLM�LIy@   $TYPES�INDEXS�$�$CLASS  ����lq�����apVERSI�ONix � ��}qIRTUALi{q'61�r5���p��q�t�+ UP0 �x�Style S�elect 	 � ���r�uReq.� /Echo��N�Ack��Initiat�p�r�
�^�m��)����	��
�� � �������������χ�q)���Option bit A<��p��B��C4�Dec;is�codY���Tryout m�j�6�Path s�egh�ntin.�8�Ig�ycX�:�T?ask OK��?��Manual o/pt.r�A����B���C� de�csn ��$�Ro�bot inte�rlo7�@�\� i�solQ�4�C��ixM�@���ment<��)�������Ě}�st�atus=�	MH Fault:����Aler�1�C�ܹp@r 1�z �j�;�y���I�; LE�_COMNT ?}�y�   Չ �ѿ�����*�<� N�`�rυϖϨϺ��� ������&�9�J�\� n߀ߒߤ߶������� ���"�����U��Ђ���Ŵ   ��EN_AB  ��:� �����������ꮵ�MENU\��y��N�AME ?%��(%$*R�זb��P� ��t������������� ��+O:s^p ������  $6HZ�~� ������/ / Y/D/}/h/�/�/�/�/ �/�/�/?
?C?.?@? R?d?v?�?�?�?�?�? �?�?OM