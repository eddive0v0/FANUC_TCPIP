��   ��A��*SYST�EM*��V8.3�0340 11�/9/2020 A   ������DMR_S�HFERR_T �  $O�FFSET  � 	  /GR�P:� $�MA��R_DON�E  $OT�_MINUSJ � 	sPLzdC�OUNJ$REF,j�PO{���I$BCKLSH�_SIG�EA�CHMSTj�SsPC�
�MOVn �~ADAPT_I�NERJ FR�ICCOL_Pz,MGRAV��� HISID�SPk�HIFT�_7 O �N\m�MCH� S��ARM_PARA�O dcANG�o y2�CLD�E7�CALIB�Dn$GEA�R�2� RING,��<$]_d��REL3� 1� N �FMSV�� +� M_LIF	��h(t*����(DSTBl+_0z*_��=�f#�&~WCL_TIM
#�PCCOM��F�B� M� �MAL�_�ECI�P�:!�%X{ g$PS� �TI���35�"L $DT�Yk9�f1END�m4�`1�ACT1T_4�22�93�94�9�5�96�6_OVR�6� GA�7�2�7�2��7�2�7�2�7�2�8F�RMZ�6DED=X�6CURLNHS�2sF�1�G�1�G��1�G�1�G�1�CNA�]1?(B0�$M��sPL� W ���STA:#TRQ_�M��k@KNVSUXZYZZYI)Z�I7ZIET �VC�MRPRU : � �B_V�:!�RHEP�TSI�Zn�SDATn �JOI���T ��T��V��X�^��9P�(ORGlNEWl��T��T��V��U� �Ys  ��$�1SS> �S���a�����`�VERSI� �g�  ��~�aIRTUAL�oܫaS 1�h� ���N  ��
C.gN� v���v�`���}�}��a��|��Ҿ �Fv��6����� =6b �g�S���q�@��������ˏG������*�<�'�`���d�P���������=L̙͸�ߟ?�����@� �%�7�I�[�m���������ǯٯ�>� ��e�$��D��d  2x�u���������@Ͽ������<d� A�S�e�wωϛϭϿπ����������`5�( N�;�J�_�J߃�nߧ� �ߤ��������%��I�4�Y���$S$ �1�lDj�S �tL�LJM���Wt�F��5U��^�@hL�F�g�D3x��;��7�;�.�(<����]� +�=�(�a�L�����
� l�����s� ��$HZ 揀eF���	�Ze�0ZrE�C�, >P!���i ���/�(/:/L/ //�/�/�/e/�/�/ �/ ?�/$?6?H??? ~?�?�?a?�?�?�?�? �? O2ODOOOzO�O �O]O�O�O�O�O�O_ ._@_�O_v_�_�_Y_ �_�_�_�_"Ҹ_o/o Ao�_eowo�o�oZo�o �o�o�o�o+=�o as��V�������'�9�b,(�$1234567890]�o��[��� ��������ُ��� �!�3�g�W�s�{��� ����͟՟���'� /�K�u�e��������� ��������M�=��Y�a�s������!(�XϿհ��PLCL������� D??�  �+��N�?r�]� �ρϺϥϷ���������8��VCMRPMR��2���dL�� ��0+ߩ߻� �ߔ��ߔ�	�#�-�� =�c�N���������