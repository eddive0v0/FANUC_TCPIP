��  �A��*SYST�EM*��V8.3�0340 11�/9/2020 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  �  �ALRM_�RECOV� � � ALM"EN5B��&ON&! �MDG/ 0 �$DEBUG1PAI"dR$3AO� �TYPE �9!_�IF� ` �$ENABL@�$L� P d�#Uژ%Kx!MA�$iLI"�
� OG��f �%CAUSOd�!PPINFOE�Q/ �L A� �!�%/ H� �'�)EQU�IP 20N�AMr �72_O�VR�$VER�SI3 ��!COU�PLED� $�!PP_� CES)0s!o81s!Z3> ��! � $�SOFT�T_I�D{2TOTAL_�EQs $�0�0N�O�2U SPI_I�NDE]�5X{2S�CREEN_84no2SIGU0o?|�;�0PK_FI� �	$THKY�-GPANE�4 ~� DUMMY1d�TDd!_E4\A!R��!R�	 � �$TIT�!$I��N �Dd�Dd �DTs@�D5�F6�F7�F8�F9�G0�G�GZA��E�GrA�E�G1�G1
�G1�G1�G �@!�SBN_CF>"
� 8F CNV_J� ; �"�!_CMN�T�$FLAGyS]�CHEC��8 � ELLSET�UP � $�HOC0IO@� }%�SMACRO�ROREPR�X� D+`�0��R{�UHM�P�MN�B�! UT�OBACKU��0 �)DE7VIC�CTI:0�A� �0�#�/`B�S�$INTERVA�LO#ISP_UN9I�o`_DO^f7��iFR_F�0AI�NA���1+c�C�_WA�d'a�jOF�F__0N�DEL��hL� _aAqQbc?Yap.C?�Y`�A-E��#%sATB��d��AW{pT $DB� g"� =S�$MO�0B x!kq� \� ;VE~a$FN!�p�d�_�t�rdTM�P1_F�u2�w1�_~c�r~b MO<� �cE D [�mp�a���REV��BIL0�!XI�� �R  �� OD�PT�$NOnPM��I�b�/"_�� m�蘁H��0DpS �p E RD_E�L�cq$FSSB�n&$CHKBD_YS�r�aAG G�"$SLOT_�H�2��� Vt�%��x�3 +a_EDIm   � �"���PS�`84%$�EP�1�1$OP��0�2qc�_OK8ʂ� e0P_C� c��+dR�U �PLACI4!�Q���( �a�p9M� <0$D������0pB�UOgB,�IG�ALLOW� �(K�"82�0VAaR��@�2�sBL�0;OU7� ,yq�`�7��PS�`�0M_Ox]d���CF��7 X0GR`0�z�M]qNFLI�<���0UIRE��$ށwITCH�sAX�_N�PSs"CF_�LIM�t=�SPEED�!���P��p�PJdV���u�u�3z`�P6��ELBOF� �W��W�pH� ���3P�� FB ���1��r1���G� �� WARNM�`d܁�P����NST� CORz-PbFLTR۵/TRAT�PT `� $ACCQa�N �r�pI�o"���RT�P_S�r C�HG@I�Z�T(���1�IE�T�Y1�݀�� x pi#�Qʂ�HDRBQJ; #C��2��3��U4��5��6��7��U8��9s!k�M$��	3 @F TR�Q��$�V����C�FN�_U�pY�k�OpT <F �������#�I2q�LLEC7�>"MULTI�b�"��A!cj DET_��R  4F S�TY�"b�=*�)�2��o���pT �|� �&$L�>�+�0�P��u�!TO���E`�EXT�יၑ8B���"2����
�t k0F�RLƯ�r�q���� !D" �M��Qm� �蠋c������"��G�1�ց�qM���P��! �����# L0	����P �pA��$JO�B,�ǰR�0�TRIG��$ d������ �� �K� l��弧�qC`�0b% t���F� CNG0A�qBA� ��x��
�!v@��� ��z�0�P{`X�R·&ΰf��Pt�a�!��"J!�_)R��rCJ$�*(J)�D�%CHӽ��z@h�P�Z�@ '.�RO`�&�ס�IT�c�NOM_�`���Sj��pTE(�@�݉��P�ǭ��RA�0�2&"<�>�
$TFV w�MD3�T���`U(C1[�g�'�Hgb�s1q*E���\Ѕs�q�ŦgAŦsA�YNTt�q�P|pDEF�!)��G�PU8/@������AX��Ģ�ewTAI~cBUFņ��|psQ* � l�'�PI�)�P\7M[8Mh9� k6}F\7SIMQS)@�KEE�3PAT�Ѡ"�%"�"$#�"�L�64FIXsQ+ �ԭ�AdC_v�����23�CCIh��5PsCH�P�2ADD�6�,AE,AG,A!H�_�0�0_,@�foA)� ԀzFK� '�=$#�"�:�4E��, l���7@zpF�CE�C!F+H�S�EDIS�G�3�-z�P��MARG����r%�FAC
��rSLEW<���x;�,M��MCY.����pJB����
aC�W�v��U��W/ ��?�CHNS_EMP��$GE g݀!_} ����pP�|!TC9f��y#a���Nd�W#%I��r<��<�J�R�И�SEGFRfoPIOj�ST`�gLIN׃�cPV����!�$0�����b�'��b�B��1` +`��	��a	`�� �a�Pܠ��At��Py�Q�SIZ���ltKvT`VsE pz�y�aRS%� ��uc@Q{k�|�`�xZ``Ld�| `�vCRCɥ��!����t�`%�p9a˭9b��MINQ��9a7��q�D�YCk�Cz��le��50�Lp ��EV���Fˁ_leF��N����Q(۶�X%+4,��#{0|!VSCA�} AY��c1G"�2 �>�
/Ψ`_rU@� +�w][��i %�7�P}R��3� �ߠ�߱���5ġR�HwANC��$LG��l�*1$�0ND�סAR�0NK�a�q��acm�ME�1��n��A0h�RA��m�AZ�����X%O`�FCAT���7`�vS�P.
ADI�O��� u��pWP ������ⁱGv�BMP�d�p�D&ah�AES�f@̓�W_P�BA�Sk�s��4  ��I�T�CSXh@�w�5��	$�K1�T��?sCb��Ny`�aBP_HEIsGH71��WID�06�aVT�AC��u��!AQP0� �\�EXqP+�L�@��CU�0_MMENU��6��TIT�1	�%���a�!A1ERRL���7 \���q��sOR�D��_IDG�=�QUN_Od�L $SYS���4��j��Iϡ	�EVG#|�a��BPXWO��z��8��$SK��*2 ��T(�TRLn��9 �� AC`��u䈠IND� DJ$�4 _Z�*1K�*��W�PL�A�RWA�.�tТSD�A�ת!��r@Y�UMMY9�ª�10���¾���:	�A1PR�q �
��POSr��;� ��[$)$�q�PL��<�ߪS�@��=�'�C�>\4�'�ENE�@T{��?S�S��REC�OR.�@H z�O�@;$L��<$��62����`_q̸b��_D9�W0ROx@�aT[���b�.�`F��������PAc�|��bETURN�V�MR��U� ��C�R��EWM�bmAG�NAL� 72$LAx�e��=$P��>$P٠= ?�y�A<�C���@�D�O�`����:���G�O_AW ��MO�a)�o���CSS_CNSTCY�@A L� ^�C`' SID[^�2
2�N��O���ـI>�� B PNP�RB^rzCPIP=OvI_BY�R}�T�r��HNDG.�C H�DQk�SP�s*�SBLIO��F��0��LSD��0N0�	FB��FE��C4��жE�DO&a-sO�MC`{�4��C�rH��WFPB�����SLA�P�F�bIN� �N3������G� $$ ���P]��v��v�ޕ����!o�"��#I!D�&L�&W�";$gNTV*3"VE 4��SKI��as�3�'2�b&aJ�&aM��mdSAFE,d�'_�SV��EXCLUt7ѻ���ONL`��#YcL���4��I�_V8���PPLY�y�R��H[0'3_�M@�NPVRFYI_S�2MS�O@���k6�1�~3�#O�t !5LS�E��35H�£1�`%�P���$��t5�%� Hy��TA2�DP���  �_SG�� I � 
$CURB�_�
�B �������#H��3F��UNM��DZD@���l�{IxA��J��F�EF��IM�J� @F]Bk��pOTb�k�ԋѭ5�׿P��и@M� NI��K���
RwPA!(TD{AY��LOADj��R�ӵ2 �EFV/�XILy��q�}�OhPe�D�_RT;RQ�QM DF�����P�r�S`�ThU 2L�`���Qk�P8���Q�QN 0�A�QaA�t�R���DUb���"�CAB�aO��B�NS�QW`ID��`PW���U/q� V�jV_�P�P���D�IAG�1�aP�O 1$Vb�HuTl�@�u�t� �j���rRp�lDQ�tVE��Y@SW�ad�p7`q��U2�PM�p�QOH�U�Q3PP�`�sIR���rB��Fb�S��q��q�@ 3r��-x ��-uj#e��PO��P���uRQ�DWuMS���uA��u�b�tLIFE Z��C�p���rN�q�r��uxA�s�rI�xBCVp���NC�Y���r�FLAW�y@OV����vHE'ArSU'PPO2���rS�1_E�)E�_Xf�h���s�Zp�Wp�p�s�0��xA���XZ����VqY2ˈC
�T��D���eN됕exAJ�% v_��q��/�Q `[ CACsHE��3�SIZ�v�*��"j�N� UFFIo� �p����$�3��6���M�����R 8�@KEYI7MAG*�TM�ᄣ���D��q�`��O�CVIE�`�S ����Ll$@)#?G� 	��%���T�Pm�ST� !� �`!��@!�VP!��0!�EMAILy�1Q|��� _FAUL���U� �9��COU�z ��T��|aV<' $��zS�PC`;IT�#BUFF�)!PF�Oy�o�D�B���nC($����Ú�SAV�Ţ�`���`���|FP
�z���d�� _���"P_�OT�����P[0�Ѓ� B��AX��-�I���Wc�7�_G�s��YN_$q'�W�RDuY��U#rMb�T���F+�fP^@D�&�X�������g�C_��&�K��8�4B3���R��2�q��DSPl���PCy�IM� pÖ��#�Æ`UM�:���K0d�IPm#�q	�o�TH��=c�mPyT��p�HSDImƏABSCz$��o�V�� �Я�&�`ӀQNV�!GO�&ԑ�mƸ�	F�aаdR����,��SCxbk(�MER|4�FBCMP3��ET�1�Y��FUX�DU���\���%2CDf���z�u��R_NOAUT�  Z�P4 �"U��IUPS�C	@�C�1ϱ	A㍰���[H *�L  t�3���֚@�0�# �����A��VQ��1��扑��7��8��9P���p���1��1��U1��1��1��1��U1��1 �2�2�몥�2��2��2��2���2��2��2 �3J�3��3���3�ꨴ2����3��3��3j �4�_�XT�aQ\ <���I�簉���3刡FD�Rxd]T��V��0���r��rRE�M�`F��rOVM�I�>AGTROVfGDT�gMXv�ING�fuaIN�D��r
��а$DG��:sp��ur�aD�VpRIV�м�rGEARI�I%O�eK7�tN�%(�hQ�x0h `��sZ_�MCMÀ�q;�U�R��^ ,�1?g �� ?� .�a?�!E�0�!!�����_P}p5P���`RI�դ$��aUP2_ ` VPģTD���3�#�?@�!�'�%@�#BACܲa T�ŢڠZ�A);@OG.5%�C8T����IFIq����x�:pC5PTV��MR2
b� �3LI ��3#/5/G/^|���u7_���R_��A�԰`M�/-D�GCLFuDGDMY_HLD�!�5�vP��tz3�c�P�9? T�FS]��d P� �B�0��а$EX_�A�H�A�1kPl���@3[5�V�G:�
e �����SW�O�vD�EBUG4WR�eG�R� �U��BKUv��O1a� pPO�P�YoP��BUoP�MS�0OO���QSM�0E����� _E f �`|Ȱ�TERM�Uyg�U���ORIe0��Qh�Ul��SM_�80Ţ�Pi�U� �T�Aij�VDX�U}P�k� -���f$�Ua`g$�SEGfjx@ELT}OV�$USE��NFI"��bn �q�+�d]dh$UFR�02���a���	@OT�gU�TA ��cwNST`PAT��<?��bPTHJ ����E�:��АbART�+��e|�+�V��aREyL<z9�SHFT�¸�a q.x_SHI�M�^���f $`�xj�)A�0OVR��ǲSSHI_p&DU4� %��AYLO��AֱI��ѻ# qk�%�k�ERV���q�yz��g`�<r4_0&���_0RC<�!9�ASYM	�9�F�aWJ�g��E�#*qV���aUz�`ֱ.u|���DuP���pYі�vOR`M�3Z�G	R�Q1Tl�oR�V�`�`A��B��m �t>�b671TOC�a1�QT!k�OPZ2��P�}���303OY�ߠREM�Rm�9�OXѐ$�reT�R�e�h�Fq/4e$PW�R�IM���rR_C�#tVIS`sb�3UD�#fsSVW�B��b n� $H|.56�_ADDR�H�QGr2�'� �
�qR��~�o H� S��Q�4_���_���_���SE�A�H�S��MN�Ap T���_����OL���v���ּP�ACRO���aS�ND_C����qٔZ�OROUP���_X���@��1��25� ��?�4 ?�<@���?����?���2AC�I	O��W�D:���J����1Sq $� ;�_�D� �PM���PRM�_.�^�HTTPu_�HQar (��OBJE��"�/4-$�LE�c���s � ���AKB_�T�SS�S�� �DBGLV��K�RLÙHITCOmU�BG��LOF�R�TEM�ī�x�e�a7f�SSQ ��J�QUERY_FLA���HW��aQaetZ���F�PUR�IO�h����u��у�ѿ� �IO�LN2u��
@Cޞ�$SL�2$�INPUT_�1�$��i�P m�D�S	L��Qav��gߢԝ�h=�s�=�_�IOయF_AS�Bw%0�$L:0'�:1�q��U`|p�aTժ�_��p�HY� ���`��U;OP�Ex `��>�����hᣐP��Ã�^����x�q�� UJ	y � �� NE�wJOGܾg��DIS�3J7����J8��7!PI��a���7_LAB��a3������APHMI� Q��9�D�@�J7J�� �@_K�EY� �K^�LMONQaz� �$XR����WATCH_� �s98.��ELD.5y� n�&�E{ ��aV�(���CTR@s����%Rv� LG�|����DSLG_SIZM�� &�@%��%FD0I$;�Q2 #�P=/" _�+� �@��ЩR ��P���S��� �ťV" ZOIPDU�r��N��
3R}J���@P�A�҈]�d0U�-�L�6,DAUREA`��/�h^GH0�}��OGBOO2�~� C��ӐI�T�Ü>@��REC��SCRN����Dx��FR'�MARG�2 Ҡ�����N�"����	S3���W���A���JGMG'MNCHL����FNd�J&Kp'7PRGn)UF|(�pn|(FWD|(HL�)STP|*V|(e0|(,�|(RS�)H�+��C�t�#y���1P#'G9U籐$"'�r0&��d�"G`)WpPO�7��*��#M07FOC�wP(EX��TUIn%I�  #�2,#C 8#Cl p!�p��v3@����p�N�sANqA�҉b�pVAI��CLEAR�vDCS_HI\T�Bu�j�BO�HO�GSI�Gr�HS�H(IGN; ���Mm!��T٤�@DE�(4LL\�C���SBU�PR`���pmT4B$1EM�נ���rRQa����pW��Ρ4�OS1*zU2zU3zQYT�AR`� ����΁�e sԲs�J`�P�r��aO�P��a�VST?��RiY��a �$EfCkW���&f9f!�U��V�� L���_�#�|p��U����וE��֕YU�_ � �� .�x6���c �MC �� ���CLD�P?�J�TRQLI��[����i�dFLG ���`��srAD��w���LDutuORG��!21r��vyxu�p�t���dд� ���`t"5�du� PT�`贴bp�t�vRCLMC�t}��y��YPsMI����� d)ֺQRQ����DS3TBP��P [���h�AX�bi�k���E�XCESy�;�M���U���`O��dE�;��V����]�_�AW�\��������`K�B� \�����$�MB��LI�I�R�EQUIRE�cM�ON�
�a�DEBU���;�L�`MA� �ڰ ᛐ����qV;�ND>S��'���ړDC�2:I9N�7RSM������@N���F3��PS}T� � 4}�7LOC�VRI���U;EX\�ANG�RY�^;�ODAQA�K�c$t�1RBMF�� ]���Y�b0�eǥ�C�SUP�e�QFX�S�IGG� � ����b�wÓc:6�d���%c�?���?�.���DATACWk�E��E������N"R� t��MD
��I�)���@��-���Hp��ᥴX�!�ANSW!��`Q�1
��D��)|��� ���� ÀCU; V0� px���LOj������5�W�3�E����U�M�;�RR2>B��� (E�N�A�q d$CA�LIa��GvA��2�9�RIN� ��<$R��SW0���)��ABC��D_J2�SEu�Y���_J3:��
��1SP���Y�P���3�"��
Y�J�J�CZ՞r��O!QIM��(�CS�KPz��1oC��Jq(�Q�ܺՠպհ׎e�_AZ�rV���E�LQU��OCMP0s�)����RT���G�1���5��P1��9�f�G�ZE�SMG00}��Օ`ER���Å�PA �S(���D�I�)�JG�`SC�L����VEL�aIqN�b@��_BL�@Y����Z�J���������YPIN�ACcR���	"x��f`_u�!�<���<�b܂�F���YPDH��t;����iP$V����'A$d�b�ȏP`��qy�B��H �$BEL��||�_ACCE��� �����IRCi_����ppNT�Q��S$PS���bL  ��&s�	1<w@
PATH��_D��_3..���_wQ �� ��rb�CC ���_MG !$DD���`�FWE�~���������DE�P�PABN6ROTSPEE�{Q�`��{QDEFb���. ?$USE_��BC%P��C�0BCY��Z�q s�YNA�A�p}yм�}MOU�NGRR� O��Q�INC�m���h�x���i�ENCS���d�Y�&��f�# IN��RI.%���NT�����NT23_Ux��`�A#LOWL�AA~0��`�a&Da0@Y�C���`���C,��(&MOS�@�MO��ǀ�wPERCH[  ~#OV�� �' �Q�#F�d"&�F��
�gm �@w�A. 5L ADw��v�)%�d*_6�z&TRK���QAY I�3쁏1.�5�3n�p�����PMOM B�h��sp"�W����0�3azR��DUЋ�S_BCKLSH_C.!E��&� ��-�?D�JJ���CLALBP'"�q�0܀|E�CHK�`�US�RTYJ�N����T:Seqr}�_c�$_UM����IC�C����C(LMT�_Lwp� T̱WE]&P[P !U,�5A�+0gT8PC�!8H�`|��2�EC�p�bXT���CN_��N���V�SF���)Vg�a	'�|�Q.
e�XCAT�NSH������eq�
A
&F�/F�Z� P�A�D�_P�E�3_ �`���6� �a�3�d�E�JG�p���cO OG|�W��TORQUY /Ւ#�9� ?��"��� r_W�5�4C��<tP��;u��;uIC{IQ{I��F��.qaҐxp�� VC��0b�Z��r�1�~���s��uJRaK�|�r�v�DB���M���M�_DL��:2GRVBt;���;����H_L��b �i�COSv��v�LN�p�������d�@��mq׊Ō�q�Z����&�MY�����T�H��6�THET0j%NK23��`��㶣�CBe�CB��C��AS���mt���󌘑e�SB��p�GTS��(C�m�=���cM��ԃ$DU��@C7����� ���Q�F�s�$NE��ؠI@���C)���T�AX������h�s�s�LPHv�_�9%_�S�ңŅ ңԅ_��������EV��V����VʪUV׫V�V�V�V�V�H��E�²P��?aٸ׫H�H�UH�H�H�O���O��ONɹ�OʪO�׫O�O�O�O
�O�F_�����Ņ��Ė�SPBALAgNCEQԃQLE͐H_X�SP�9��ņ9�ԆPFULC�=�d�L�d�ԅ&�1���UTO_�@�eTg1T2����2N�A ��?�Ԗ��1f�D�5���1TP0O����,p�INSEG��!R�EV�փ "!DIF�y5K�1�0��1��l0OB&�lAE��72�p?�A$�LCHW3AR��AB�a�5?$MECH��%�X���FAX�1PJTp��z���З 
��q�%ROB� C�R.��R|���MSK_���� WP ��_WR���r0�?{41	b4 2`0�1#JD0���IN���MTCOM_�C�p��  �� 8�$NOR�E$#���t����� 4�0GRr��F�LA�$XYZ�_DA��TC DE�BU�� ��t��u 0�$uCOD[AG ���2���0�$BUFIND�X2 ��MOR#�� H-��0����FB �0�JD$���c�QVPTAA�+�2G6� �� $SIMU�L�` 13�3O�BJE;ТADJ�US�� AY_It�A	8D�OUT�`����0�_FI�=@T+p4 ��X�3p3�A�5DNrFRI(CXT8E�RO�` E3q[0��OPWO�p'�}, SYSBUq�( $SOP��A�U�3�PRUN,v��PAC�D��℟0_� NR�X�A�B��PP� IMAG�[A-�G�P�IM�Y"$IN,��!#RGOVRDM�� ��P   #`W�L_`��an%�B�PRB5P�X�`QMC_EDT/ �� PPNq�M�"<OQ@MY19NQ+ �M!SL;�'� x $OVSL��wSDI{DEX�S��&�SP1�"V3p�%N 1q�0378�"zA�$_SETp'� @�0K2��AASRI�� 
^6_��j7�1v1!+ 5� �P� �<T���`A�TUS@$TR�CI�H%�3BTM$�7�1I��$4NQ�3\� '� D-�E��"�2z�Ev��1!0l@�1EXE�0�A�!B*B�4S3�Z0.��03UP��9A$Y�' XNN�7�q�$�q�9� �PG���? $SUB�1����1�1�3JMPWAeI,`P	3�ELOP����$RCV?FAIL_CH��AR-���Q�P�Tx�U�R_PL�3�DBTB�a�R�B3WDV��UM�`T�IG�( ��4`TNL(`TjRRm���`$
p	1XQ� E�S�T|�R�ADEFSP�� � L-���Pq_�P��SUNI#��7�PmAR1@��3�_�L�P�1+ Pw�&����`�� "<0���)�T"NU�KET(b(p��`P^R&��� h� ARSI�ZE� ��1��naS�� OR�3FORM3AT��TTCO� ja��EM���d�SU�X�2l`�PLI�OR&�  $>��P_SWIu��!��fLLB&�?� $BA�`1�3ON9AKPAM�0=<y��BAJ5����2r68v��_KNO�W8cNrA�U9AߐD�x� �PDC�ryPAY�[�t���y��w�Z�sL�1��U!PL�CL_$� !� �s,qv�tb"z�vF�yCRPO�zL�2�tES���wR4�x�w�tBASE$�J��W�_J�qK�mA��fBu��r�q�"+ MAX4P�`AL_ � $�QPh 1q�!��C[�D�s�Efr�J3�����{ T� PDCK� |��T"CO_J3�������
�hr���� �桀C_YQ�  �s ��ЏD_1�z2�tD���n�^����m�|TIA4��5:��6[�MOMS ���ȓ��ȓ��B�@A�D��억��PUB{R͔������e#��` I$PI�$�QM�=q�w k�B1�yk���������iqRM�q�!Ħ~AĦA
��9d5SPEED�G�b��E �T��T�EP-�C���Q+�Q�ESAM (�E�����Ep{� m�$�� k� ��~@Ƕ�P_�ֹm�k�@v{��ŵ��,H��ǳIN̚�c��1ˀ��B�W�.�W�w�G�AMM��1��$GGET9" �D;�zu
��LIBRcA��RI��$HIb@_�=!�0k���Eh ��A����LW��4�+܀�X��7���wP��C�EUv�[ �0 �I_b�xu��L� ������ȓu��ٞ�� �$Ј �1���I�0R��D`\��kAT��LEf�=q�1M�7�ୄPM�SWFLTM��SCRsH7�����!���~B�dSV&�P�� A �����#S_�SAqs$��eCNO;�C�1fB<�����K� ����S�C���hrǥ��m�D� a���� �� �в����U!C�p�������s �c}MJ�� � �ӣYLi�K���^S J�|v!6O�K���@BK�- ��OW����9���M $P��p����Dc�"���1~B�`M��T2�� � $-�$s$W� �%ANG" �q� ����!�� 5P&��o����c�#J��X`O"���Zz��`�@� �y�OM��+�(�:�L�^��p���CON@�U Jt�b;�_�B� |� ���ș@&��@&�����m'X&��.��� 9�'�� �`"&�Pma�PM0QU��� � 8#`Q�COU���QTH�YPHO/� HYSf�`ES-r� UE� ���S`O�d�   �$P�@�Ŋ2UN��0b�@O��  � P�p45�E��C�R�ROGRA�1A22DO445IT�Ё1�F0INFO�� �%0g;�1AȬ!O�I�2� (�SLEQ���1��0k6E1yS�НD� 4#`�ENAB"20PTION�C�T̢/G�T�CGCFA� @b#`J$P��<2����RdH0OBG�2S�_ED�@  � ��{K�q�3��E�)�NU�G�HAUT<�ECOPY�qI0(�L���M��N�@�K^��PRUT �B�NV@OU�b$G�92DT�!RGAD5J��bbX_ �RC$`pV�pVWnX�PnX[�pV�`Pz�N^��_CYC"ZS�NSE�$ ��LG�O���NYQ_FREQ0�Wb��a�d23L�p�b�PnQÓb��5CRE���#�гIF��s3NA���%?d_G��STA�TU' ��*7MAI�L��YsIN��$LA�ST�a���TELE�MA� �GFEASIA���� H �b�1���f;B����I�0���R=q�!� R�&rAB+A��Ex0��V�a7vW�Cy��1�U�8�I0�pd�lvRMS_TRs��@� �sr7�z��aktB�R��/ 	�b 2� =�_+��v e��w�r� �fe���c�G�DOUa3;�NLHC�RPR	 @��2�GRID�1+CBA�RS��TYC�RO�TO㐾�³�&0_"[d!�P��B�OxD�� � �0�P�ORa3��[���SReV_`)˄ÆDI�T^���������U4��5��6��7��I8ぬ!F��A�#0?$VALURs����d�q_�D�� !E��u1��aa��F=@AN�㉒qaR�@|a��TOTAL��,1��PW�SIJ���REGEN����#�XxxI3e%!��� T1R^s0���_S��^���CVnQ�D��B8rE�cN��!��42�@Ó7V_Hk�DA�~����S_Y
�rfS���AR�2� ><RIG_SE�ch�dÂ�e_80��C_v�~`�ENHANC�!O� p�qEqb�ý�INT��� yF.3MASK��.ipOVRFcP� N���`a
�_�*6^�M���B[��f8��SLG|����� \ �� eH ���Sq�dDE�U��*7Ő�d%��U�!�TEj>  � (7���↡J϶�"cIL_�M!d��P㈠�TQ@� �Ë1rpj�eV�ˍC��P_��op��M���V1��V1��2��2��3�3��4�4���ᄠ�����؃�s��IN��VIAB� �İ����2��U2��3��3��4��4�ؾ���#"��������%��׌ՠՌ�PL�v`TOR� ��IN�b�����  �p���MC_F� 	����L����B�ڐMb�IB���#� 1 ��)���KEEP�_HNADD��!H��<p��C�_`������H ��O�!��P�������G���REM���쑥�;�R�W��U[de��HPWD�  ��SBMTo���G�1�2��� H COLLAB u��a������ؑEb�0IT���0��n� ,� FL>bq$SYN���M�C��d�UP�_DLY��#2DGELAJ �nbY� �AD�� QSwKIP�� Ļ��60ODD���t P_ 60_2�g0^ ��� �		Q�	��	%��
2���
?��
L��
Y��
9��Q�J2R�P�ΊCX]pT�SY���X]P��Y�1�� RsDC��b�� ��@	ReCg�R4ae��"d���RGEr@sl�:��FLG�!Pa�SW��I��SPC�3�QU�M_Yt�2TH2�N&�# L 1�� �EF�@11�!� l�����C��AT4�ET1� �7s"k0o4j!�@Y�j!<<3\�HOME�"�P
<$2D"�J/\/n/�/(�/�/�'3D"��/�/��/�/?!?�'4D"ӀD?V?h?z?�?�?�'5D"��?�?�?�?	OO
�'6D"�>OPObOtO(�O�O�'7D"ֻO�O��O�O__�'8D"׀8_J_\_n_�_�_�%S��1�9 �q=#$����S�E���·��LbݖJcIO�q�jiI�P���GbP�OWE��� �4` wGbה y��b$DSB�GGNABqՔE C) z���S232Pe'� ���U�P�OICEUQrt�E3 >��PARITáՑ�OPB��FLOW�TR`�c�3�ֶ�CU+pM��UX�Tn���U�ERFA�CtC�Uѐv�bCH�q� t��b��_p��$�����OM۠9�A�T\>���UPD�A#�`T+`҃*�� �x�s!��FA�������RSPqpQ���� !�X$USA� ���Y�EXmpI�O6��pU�YE��b_`�ª�B�#q`�WRp���_�YD�����VF�RIEND���U�FRAMδ��TO;OLȆMYH�����LENGTH_V�TE��I���[��$SE�`��UFI�NV_�@�5aR�GI���ITIĳ��XX�	�J�G2J�G1T�U�D�d�u�2��_Â#O_p�p y�ၻ��n�C	�z��C ���ʖ ��G��zr2�� @ 9�qC���d�wu���ysF� ���p���X #�E_M�pCT^�H��f��(<u6�	�G#WV�z��G���Dh LOCK~�U� ������{$� 2���H~�D ��1���2��2�3��3���:� ���V��V=�"�=�F��V��!Ѕ�/�(⑪��p�xṿ ����Prƻ���������E������!�6�AC�PRs�D!�}�S���`���<��a� 0 5�"ؠ�V��ؠ���	�������
M�S��� ح�R�qda�¿$RUNN�`A)X2q��A��L�+"^��THICx� �w �u��FEREN�g���IF��x���I0����V��G1&�*�Є�1ٲ[�I�_J�FR�PR��
��R�V_DATA�q� RD�[ 
�A�L� �xՑ ��b{�  2� ��S��`�	ܧ �$ Z"G�ROU��!TOTܸ���DSP��JO�GLIYs�E_P�PrO��\7`��bv=K�p_MIR�.�2��MQ�O�APp���E<�o��t��SYS�E�ib��PG��BRqK���v$ AXIa  �⃃���Ҽ��A����H�BSOCd��T�N���16��$SV1�DE_�OPNsSFSPDO_OVR4 ����D� �OR+��PN��P,�F��,��OV��SFa���d�$�F�}�ja2㒓��ҁibL�CHH\RECOQV�n��WE�M�����RONs���_����� @�9�VsER��n�OFS9�C�Я�WDE���A����Rh��TRBq|6aY�E_FDOh�MB_CMkS B��BL��.�u��8āV摁��p��]�Gv��AM��i ������_M� [r�ec� T$CA��D:��HBK�q�vIO��,�a��PPA L1\D���bDVC_DB<���q�b���ja"�1���3���/ATIOi`jqcp��U�� �efCAB �����J���������__p�vSUBCPU�b�Sv��`_ ��p"�`'}���b"�?$HW_C� IpȺ��'ɣAx����$/UNIT��� � ATTRI���"��CYCL��NEC�A�Y�FLTR_2_FI#��h��fƂ�LP$���_S�CT��F_�'F_�,E2�*FS�a��"CHA��-7�1�Pr�2RSD  �b������a�`_T�PROX�MFpEM	`_��r��Ts2�� s2̍��5DI&��tRAOILAC���M��#LO�����5��ﰰ�����PR�S�̑{�dAC�p	���FUNC!��RIN됫�|�@�DEq3RA�@�� �C87`�CWARB�	#BLƑ�G�DA�K�!�H�HDA��AX�C�ELD�p�@S��2�A�@STI��`U��ѓ�$<�RIA��q�bAFQ P=���S��U ����3MsOI� PDF_�ؔ��qHpLM�FA�E�HRDY]�ORGEPH�0��|� P�UMULSE���`'*���0J(�JC�X��S�FAN_ALMsLVBs_aWRNfeHARD���v����p�@2$SHADOW��0��a�b��_`�+q�ї�_���vAU��Rx4\rTO_SBR��e���j� �|�A	sMPINF����!t6Q'sREGL���aDGBP��V�pL.�l�FL�%!���DAՀ_�P�C�M��N�Y�B �8V  ��� ]����$N�$Z�� ��Ҭ����� ��|�EGK�����qAR��#��2?��wP��AXE��ROB.��RED��WD���_F���SY��!���:h�Sr�WRIE��v� STR���`��7�E�!�����a���B����@CD� O�TO7q����AR�Y����.A���#�F�I��9�$LINQK�Q���y�_����6��8�XY�Z�bB�7P�OFF�
 �7�+��B��yB�����0}@��FI� ������yB
�_J��5������`Ȅҋ8��H�T�B�b�C0x�D�U �9AETURBa`XgSW���rX���FLz���#�p�u�Y���3\��� W1��K�M����31�DB`%��`'2ORQ�6�ѳC��}� DB��>��P��%����ќ\q:�OVEA���M 90=ѻs[��s[��rZ� �`X��aY�� X�O�~@ 91�P��B�F����=� S�B�_���s����SER�A	EBE��H� QC"�Aб������E�2��Q&QAX ���Q� �!�|�A ��+a�����@@��O����n������N���1 ����`��`��`�� `��`��`��`�� `��`�!��� �R�g�DEBU�#$��A�c�2��3�AB�GE�;�V�" 
�Ҷ���z!$� 
�$��$�@A$�O�$� n�$��$�N��T#��R\����LAB���� �GRO0��l� B_�1	ƞ�>� ���`�������a	�ANDàE ��<���aF� ��q��Z�0Qi�� ;�NTq`�cR�C�1=��
��{J �pERVE��N�p� $q��@A�a!��PO�`X `�����Q�p�p�$��TRQm�
���Q�����R2��oP@_ � ql=���fERRҒ��IV����gTOQ����L%��Ď�z�0G��%%�"��|?�!P � ,��2 뺱RA� 2� d�D�pܸ  �p$`O��2�PvµOCQ�� �  YC�OUNT���FZ�N_CFG��� 4� ^v2T�d�"����m W k!E�s� ��M�08b��`���X��0�FA~P���V�XA����H��0���O A�P�b��pHELkpN�� 5ސB_B;AS�#RSR]vm@E;�S�!YQB 1��B 2e*3e*4e*5*e*6e*7e*8�5!�ROOGP� �:�NL�q)�AB��@C �ACK�INT�80�sU�``x1�)_cPUA��b�2OU��P�@^x"#�y0��b��TPFWD_KA1RlfpZRE���PqP�&Q�@QUE]z�ROB�2����`�aI b`�"#8�$C0Bv8��SEMա�6�`An�STY4SO�0�dDI1�@r�1a��Q_TM�sMANsRQAF8�END�d�$KEYSWI�TCHS3h1#A�4H}E2�BEATM�cPE�pLEks1��J�HUg3F�4h2S(D�DO_HOM�POl�a� EF"�PR�� �rS����v�@OaX �OV_M���`pP�IOCM$��7���##HK�q� �D5�_w�U�b�2M��p�44�%�FORC�csWAR�R�p!%O}M�p � @��T˓�`U��P�1�V2�V3�V4���Ox0L�R��^xU�NLO.0�ddE�D�a  �$$�CLASS `����.a�p�p �#`S�0+h�9`��?aIRTx?�,o>`AAVM���K 2 je� 0  G�55a�o�h�o.�m �l	�m�pk`��o2v7u�lV}b�ah��̷t{`BS4�� 1�Li� <��� �2�D�V� h�z�������ԏ� ��
��.�@�R�d�v� ��������П���� �*�<�N�`�r����� ����̯ޯ���&� 8�J�\�n���������@ȿڿ�����rC`�cAX�� `���s7  �%�IN.�@��$�PR�0XEQ��}�`�_UPMIl��ja{`L�PR �ji`��tLMDG ��g�`��PIOF �k`d� �0�B�T�b�߅ߗ�x�߻���, 
� ��n��o�0�B�T�g��x�������yNG?TOL  �{�p�A   ��
�{`P�d�O �� @��=�O�a�s�6b�  ��u���2b�������� ����&J4Z���������� *<N`r�~�zPPLICA�1g ?je}�����Handl�ingTool �� 
V8.3�0P/58��?
88340��sF0!�755�����7DC3x�����ޝ��FRA� ;6*-  !�� GTIVqŵ>��#AUPn1�R:b\�PAPGAPONf`�.za�� OUPLED ;1�i� /03?�E?W?�_CUREoQ 1�k  P�
a7a<�n�?�d}���33b9b �3��4H�522��:HTTHKY �?Kx�?�?ZO�?6OHO fOlO~O�O�O�O�O�O �O�OV_ _2_D_b_h_ z_�_�_�_�_�_�_�_ Roo.o@o^odovo�o �o�o�o�o�o�oN *<Z`r��� ����J��&�8� V�\�n���������ȏ ڏ�F��"�4�R�X� j�|�������ğ֟� B���0�N�T�f�x� ��������ү�>�� �,�J�P�b�t����� ����ο�:���(� F�L�^�pςϔϦϸ� ����6� ��$�B�H߀Z�l�~ߐߢ��6s5T�O��/�#DO_C�LEAN�/�$6�N�M  �� �a?�������g>D?SPDRYR=�p5HI� `�@q�8�J� \�n�������������p����m8MAX� ����17.X�-!�*2-!�"PLUGGp0�*3�%PRC��B^�b�'���O���
�SEGF� K���^�p�8�J\n���LAP�(�3���
/ /./@/R/d/v/�/�/|�/�#TOTALP|y	�#USENU�"; �8?�2s0R�GDISPMMC�� o1C�@@@$
�"4O�5 3�_STRING �1	�+
��M� S�*
�1_�ITEM1�6  n�-�?�?�?�?�?O O'O9OKO]OoO�O�O��O�O�O�O�O�O�I/O SIGN�AL�5Try�out Modeގ5Inp?PSimulated�1�OutQ\O�VERR� = �100�2In �cyclEU�1P�rog Abor�[S�1;TStat�us�3	Hear�tbeat�7M?H Faul�W�SAler�Y_ oo $o6oHoZolo~o�o�o �;�?�o �o);M_q ��������p�%�7��oWOR�  �;o��oI�������͏ ߏ���'�9�K�]� o���������ɟ۟�PO�;�Q����� 6�H�Z�l�~������� Ưد���� �2�D��V�h�z����DEV ���*���޿��� &�8�J�\�nπϒϤ� �����������"�4�PALT�m[ч� 5߃ߕߧ߹������� ��%�7�I�[�m���������I�GRI 3 �;��s���'�9�K� ]�o������������� ����#5GYk��� R�m��}� ��%7I[ m������x�/�PREG_� H �!/o/�/�/�/�/ �/�/�/�/?#?5?G?�Y?k?}?�?�?�?]��$ARG_o�D �?	����1��  w	$V	[
H�]
G�W+I�0SB�N_CONFIG� 
�;IQHR�CACII_SAV/E  ThA_B��0TCELLSE�TUP �:%�  OME_IO�]\%MOV_qH�@�O�OREP��_�:UTOBAC�K�ASMF�RA:\5+ X_5&�@'`�P5'�dX� q^ ,H5-�_�_�_�_�_*o]T���0oXojo |o�o�o�o5%Eo�o�o &8�o\n� ����S��� "�4�F��j�|�����p��ď֏��  PQ�_3S_\ATBC�KCTL.TMP� XLED.GIF _$�6�H�Z���ZrDfhD0PIN�I^��U[E-SMESSAGw@���A|�0��ODE_D�@�zFDV��O��ǟ-SPwAUS'� !��;? ((O�2� 1��Q�?�u�c����� ����������;��I����TSK  �
�d__0PUPD�T����d��ԖXWZD_ENB��WJ��STA���1��~�1WSM_CFO@��5]E�7�G�RP 2� >	BB�  A���9�XISI@UNT �2j��C � 	�z��� ��G� �Q� S�c� ŝ ���5*�����ϯ������� �4 �Ǘ '� Q����+���(�a�d�MET� 2u�PNߧ�J߼��^�SCRD�1���P�EB ��$�6�H�Z�l�~�]_5*Q{I�������� �(���L���p������������1�k��73QG�Rn����	��NA��@�;	3T_�ED��1�
 ��%-��EDT�-���J��U /��Uq4Rz5*,B�&o�Fs&  ��2�K�wʹ��E��	�-3 �X5/|�/|/��k/�4�/$/? H/��/H?�/�/7?�/5�?�/�??��?@O[?m?O�?6LO �?�O�?�uO�O'O9O�O]O7_�Oe_�O �A_�_�O_�_)_!8�_�1o��o@xo�_�_go�_9�o o�oDo��oD�o0�o3�oCRS_ ���]��Ug���	 V NO_DE�L'GE_UN�USE%IGALLOW 19	���(*SY�STEM*��	$SERV*¯�Ȁn�REGх$���ȀNUM���	��PMUt����LAY�Я��PMPAL��J�COYC10U�h�R�<V���ULSUH�
��j��ӃL��ݔB�OXORI��CU�R_ʐ	�PMC�NVD�ʐ10|~�0�T4DLIȰxß�ˋ$MRߎ�&�&�ϲ����̯�ޯ���y	 LAL_OUT k���(WD_ABO�Ro���m�ITR/_RTN�����m�?NONSTO	И��� շCE_RIAS_I������˰�F��U�c����_LIM߂2�` �  N���Nϯ�<��m�`������@ϡϳ��ϯ��
����p��PARAMGP 1U��Ύ�O�a�s�>2�C>  CV���Ef��z�ߵߗЇ��U��Ж�Р�Ъ����Ԛ٢����������C���ǀ C�j���+���?�ɲ{HEC�ONFI��w�E�G_P�1U� 49������������E�KoPAUS�19� ,�uG�Y�C� }�g������������� ��1U?e��!�M��NFO 1�(�� ��=���� Aj������}�)L��S5�!և�Ad�l� D�lzD�D�hB��*��hv��*�4#˰O�������COLLECT�_�(��pE�N`���\�IND-Ex(���!��1234567890�����$���H,��)'/L/ �|&/8/�/�{j/|/�/ �/�/�/?�/�/?e? 0?B?T?�?x?�?�?�? �?�?�?=OOO,O�O�PObOtO�O�O�"� ΀ ɶIOG "�����`O_a_s_�_WTR�K2#](�8Y
�O�^P�$,]�Z��Y�_MOR"�%� �9�Fe�Fi^oLo�o@po�o�kb�#�&-mB�?>�>����a��Kt�A�PM(<���a�-=�O as�ϗ�����^�@
����`� *c�PDB�O*���Ecpmidbg�C���U�:�  +��g)��p/���S�  �� �e�-�̏��3�j�~�1��v�L�����������g�^�)�������fM���w���@ud1:˟���Z�?DEF )o7S�)ߑc�buf.txt��M� �p�_L64FIX +�Q���˓� د��ɯ��2�D�#� h�z�Y�������Կ��ſ
��.�f�x�_E ,� �l�~�`�Ϣϴ���p�IM�C�-�]��6��>̿��=L����M%C&c.�SdF�'�
%d/5ݤ`tձv���B!!�*�B����B~��Br��BA��B�����B�-6D�B�"DaaD�C�s�D�D���D�� �FB�nF���F�E���FJ"\�y�bG��gM1�\D�y��~�}���`U�x�C�ÇЯ�д  D>w�4  E	
���Ee�3Ec���Et� F�3�E�ŚF�B���F���F�Y�fF�% G��� G	ڳH��3���  >�3�3 ;���a�v � nf��q@�a5Y���b�pA�a�t�<#�eDQ�7����F�RSMOFST� '�f�G�T1�#`DZ�2!��X�Q�;�0�R��L�?���<��M��TEST�0���Rz3SMx�-C�A�z�e����| C��B�f�C�pn���N:d�b2Iy�4<2T_�P_ROG ,k%^��/%PNUSER�  �1��K�EY_TBL  �-e1]�(��	
��� !"#�$%&'()*+�,-./�:;<=>?@ABC��GHIJKLMN�OPQRSTUV�WXYZ[\]^�_`abcdef�ghijklmn�opqrstuv�wxyz{|}~������������������������������������������������������������������������������������������������������������������������������������������A� L�CK#D#ST�ATi/0_AUT�O_DOG㺒�+INDT_ENB�/� �"��/�&T2<�/6STOP�/�"wSXC� 25K��p8
SONY? XC-56Q{���p�@����	�( АX5HR5�x-tx?�>7�?�5Aff�:�O"O �?GOYO 4O}O�OjO�O�O�O�O �O�O_1__U_g_�\�TRL� LETE�6 �)T_SCREEN -j�kcs��PU�0MMENU 1=6� <O\� o�u�_oIo��&oLo �o\ono�o�o�o�o�o �o 9"oFX �|�����#� ��Y�0�B�h���x� ��׏��������� U�,�>���b�t����� ��П	����?��(� u�L�^���������� ʯܯ)� ��8�q�H� Z���~���ݿ��ƿ� %����[�2�Dϑ�h� zϠ��ϰ����b��S_MANUAL"?ޥQDBCO� RI�G�Ws)DBG_E7RRL� 7�[��a���ߴ��� OџNUMLI I����dD
O�PXW�ORK 18����&�8�J�\�n�D�BTB_�Q 9T<����K,�DB_AWAYWӽ��GCP D=����_AL �/��BS�Y!0�UD H�_q�W 1:����0,R0��T�PA�~���_M&� IS� ��@� ���ONTIM�W�&D����
2#�MOTNEND'�"�RECORD ;1@� �����G�O�N<���� z���G��N r'9K��� ������� #/�G/�k/}/�/�/ /�/4/�/X/??1? C?�/g?�/�?�/�?�? �?�?T?	Ox?O�?QO cOuO�O�?�OO�O>O �O__)_�OM_8_F_�_�NO�?�_�_�_�<_�_�_�_'o�N��(o_oqo�_�o�o�o�o�N���o �o9$2o�O�� �&��\��5��G�Y����TOLEoRENC��B�����L��O�CSS�_CNSTCY ;2A~� h���Џޏ����&�8� J�`�n���������ȟ�ڟ����"���DEVICE 2B~� ��r������� ��ϯ����)������HNDGD C~�Cz<���_LS 2D\�;� ����Ͽ����=����PARAM �E/���?�)���SLAVE F~��J�_CFG G�/�)�dMC:�\��L%04d.'CSV(��c���6�A ��CH��n�An�)��=�[��)Ɓ-�Z�j�X�W���JPъ�C�_CR�C_OUT H��<�+ϑ�SGN� I����\��18-MA�R-25 08:�33��)05>��16:01���� Ze�7-��)�)�*���o��I�m��P�uG��=��VERSIO�N ��V�3.5.20��E�FLOGIC 1�J% 	���* ������PROG_ENB��.��ULS�� ,P����_ACCLIM^����Ö7�?WRSTJN����)��MO�
���x�INIT K�%
��) v�OP�Tp� ?	����
� 	R575�)���74��6��7R��5��12�����6����TO  ���@���V��DKEXd�d��x��?PATH ���҇A\���I�AG_GRP 2�PI�|O�	 �E7� E?h� D�� C�� C ��B�́�C��nk������C��C�m�B�N�B�zoOB�)�B�k�f3�83 6789012345���B��  A���A���A��A�O�A���A{+As��Aj�RAbJAY% x��@���p��G!��Ae�����B4�h���x�
"�����"�Q�A����A���A����A�� ��hA�x~�Ao�7A�f9X��?$>��mF/X/��h����(�"_�AY�;�AS�TAM�^�AGdZA@��A:bA3%A+�-A$����)�/�/��?�*@��;d�6���@{��@u�-@o��@i�7@c�C�@\�j@Vs{N?\0�5?b?�t?�??@_��@�Z^5@T��@�O�@IG�@�C33@<��@�6�+@/<@(�`J?\?�?�?O�8s�� nE�@h��@b�!@\�0V�ff@Pt@Ihs�@B��@;� bOtO�O�O�O�'6]^_ p_N_�_�_0_z_�_�_ �_�_$o�_�_
olo~o \o�o�o>o�o��C"��!30�2KA�@^>8�Q�r��R?��  *u^7�Ŭ�Fr'Ŭ5AF<Ru^@�p�nv�@�@�pppE�@[ A�h���uC=+�<��
=T���=�O�=���=�<���<��p�q�xG� ��?� �C�  �<(�US� 4rjr�D@����"�A@w�?f�oX� �mf����������ԏ�n��
��.�@��i?�#�
b��\>x�pn�^��G���G�^x���R�����^8�ۑ�5甮��CnB�L�]_u��&�P;�'f�d��aQ{����dD�  D� � C΍��̯ޯ �8�?Vv����>�z��
t�? ��?Z��p���C�e>����DlzhD�/Dh&x�:O�ǯPD�ïh�������3*�B��)��?h}��*�V�׿ R�����
��UϤt��gh���=��t�> �=>��ZX��m�Yϧ� CT_CONFIG Q-y��#�c�p��� STBF_TTSd�
����C�tV����MAU^�����MSW_CF���R-  _ ��O�CVIEW�SY�i����߶��� �����ߩə�.�@�R� d�v��������� �����*�<�N�`�r� ����%��������� ��8J\n�� !�����" �FXj|��/�����//j�R%CR�T�e&�!�,. V/�/z/�/�/�/�/�/��SBL_FAULT UI*n�1GPMSK��$7���TDIAG V���e�2�UD�1: 6789012345�2��?�P�Ͻ?�?�?�?OO )O;OMO_OqO�O�O�Op�O�O�O�x �>��;�
�?%_��TRECPZ?l:
z4l_?� �?�_�_�_�_�_�_o o0oBoTofoxo�o�o��o�o�o�O_/_U�MP_OPTIO1N�>*qTRR���:!9KuPME��>�Y_TEMP  È�3B���p�A�p�tUNI�7��şqF�YN_B�RK WY�)8E�MGDI_STA��u&��q�uNC�s1XY� ��o7�*�~y���d ������ Ǐُ����!�3�E� W�i�{�������ß՟ ����Xu"�4�F�X� ���f�������¯ԯ ���
��.�@�R�d� v���������п��� ���%�7�I�[�u�� �ϣϵ���������� !�3�E�W�i�{ߍߟ� ������������/� A�S�m�w����� ��������+�=�O� a�s������������� �����'9Ke�[ �������� #5GYk}� �����/ 1/C/�oy/�/�/�/ �/�/�/�/	??-??? Q?c?u?�?�?�?�?�? �?�/O)O;OMOg/ qO�O�O�O�O�O�O�O __%_7_I_[_m__ �_�_�_�_�_�_Oo !o3oEo_Oio{o�o�o �o�o�o�o�o/ ASew���� ���_��+�=�Wo I�s���������͏ߏ ���'�9�K�]�o� ��������ɟ۟�� �#�5�O�a�k�}��� ����ůׯ����� 1�C�U�g�y������� ��ӿ���	��-�?� Y�c�uχϙϫϽ��� ������)�;�M�_� q߃ߕߧ߹���E��� ��%�7�Q�[�m�� ������������� !�3�E�W�i�{����� ����������/ I�Sew���� ���+=O as������� �//'/A7/]/o/ �/�/�/�/�/�/�/�/ ?#?5?G?Y?k?}?�? �?�?�?���?OO �?K/UOgOyO�O�O�O �O�O�O�O	__-_?_ Q_c_u_�_�_�_�_�? �?�_oo)oCOMo_o qo�o�o�o�o�o�o�o %7I[m �����_��� !�;oE�W�i�{����� ��ÏՏ�����/� A�S�e�w��������� ������3�%�O� a�s���������ͯ߯ ���'�9�K�]�o� ��������џÿ��� �+�=�G�Y�k�}Ϗ� �ϳ����������� 1�C�U�g�yߋߝ߯� ɿۿ����	��5�?� Q�c�u������� ������)�;�M�_� q�������!������� -�7I[m ������� !3EWi{�� ������/%// A/S/e/w/�/�/�/�/ �/�/�/??+?=?O? a?s?�?�?�?��?�? �?O/O9OKO]OoO �O�O�O�O�O�O�O�O _#_5_G_Y_k_}_�_ �_�?�?�_�_�_�_'O 1oCoUogoyo�o�o�o �o�o�o�o	-? Qcu���_�_� ���o)�;�M�_� q���������ˏݏ� ��%�7�I�[�m�� �����ǟٟ���� !�3�E�W�i�{����� ��ïկ�����/� A�S�e�w��������� ѿ�����+�=�O� a�sυϗϩϻ����� ����'�9�K�]�o� �ߓ߭���������� �#�5�G�Y�k�}�� ������������� 1�C�U�g�y����߷� ���������-? Qcu����� ��);M_ q��������� 	/%/7/I/[/m// �/�/�/�/�/�/�/? !?3?E?W?i?{?�?� �?�?�?�?/OO/O AOSOeOwO�O�O�O�O �O�O�O__+_=_O_ a_s_�_�?�_�_�_�_ �?�_o'o9oKo]ooo �o�o�o�o�o�o�o�o #5GYk}�_� �$ENETM�ODE 1Y�U��  
�P�P�U��{�p�RROR_PRO/G %�z%�V��&��uTABLE  �{oe�w�����w�rSEV_NU�M �r  ���q���q_AU�TO_ENB  q�u�s�t_NO΁� Z�{�q���  *��������Ā+�*�<�N��HIS���Q�p��_ALM 1[.�{ ��T��P+O�˟ݟ����%�S�_����  ³{��rj��pTC�P_VER !�z!�5�$EXTLOG_REQk�s�ቼ�SIZů���STK�������TOL  ��QDzs��A ��_BWDJ��؆�K�ԧ_DI9� \�U��t�Q�rU�STEPa�s��p>��OP_DO��q�FACTORY_�TUNk�d̹DR_GRP 1]�yށd 	e�#��p��x����� �n��So �k� ���W��i�z���A���B����B�ƿBF���B-G*A�G�*ͥQ@�BK1zϭ����������<�'�`߫�>���Z@���?����>�քj�
? F�5U������ѓijߢ�V߈��E7� E?p gD���߄�D�%���  C��߃�B��  ;�  Ay@E��@UUUc��UUo�&�>�]��>П��޻� =E�F@ �ѿ���L���M���Jk�K�v��H�,�Hk�=�?�  �Q��9tQv+�8����6h�%7�����Ҿ Fv���6���� =6b �g,��FEATURE �^�UK��q�Handlin�gTool �� �roduCh�inese Di�ctionary���LOAD4�D St��ard���  NDIF�Analog �I/O��  d �- ��gle S�hift��F O�R��uto So�ftware U�pdate   �J70 mati�c BackupΦ�art Hgr�ound Ediyt���708\��_amera��F���D pr��nrR�ndImM��PC�VL��ommon� calib U}I q.pc��nf� Monit{or��wset��tr��Relia�b	 ��jp D�ata Acqu�is����� DiagnosD������ Docume�nt Viewe����
PC u�al Check Safety�� act.E�nhanced �UsGFrw ��\�weqpxt. oDIO � fi+� t\j7�en]dxErr� L*�  � �{s  $��r�� :����T "� FCTN_ Menu`v���t I�TP �In�fac% � 48\� G_ p� Mask Ex�ctg�� o��T� Proxy S�vH  5p��i�gh-SpexS�ki� " #1���#�mmuni�cC ons�apd�!ur ������"connecwt 2Pdin� �ncr stru�� I KAR�EL Cmd. �LE uaG"t\i�a�%Run-TiN�Env��"K��el +G sE S�/W�Li�cen��[GER�  �Book(System)��� R5� MACR�Os,x"/Offl� �Pa� MH��- �: \ac�1M�R� �)��Mec_hStopV!t�  ��0i���Mixx��E ��
� �0od
 wit;ch��Loa� �4z.�6 k G�1�3OptmUHM GGNW filG� HFz��g�' pmfO Multi-T= �i�4pa�PCM� fun�'{3M"PQo[�D QV�H�Regit0r�  � mpo� Priz@F�K _fcs �W g Num S�el�5��� DS� Adju� ���`W�
 4 S|Xtat�uQ/bUC�� �RDM Rob�ot��scove��� cctO Re�m�0�n���SS�ervH10@#CTX�PSNPX yb<2�� "K9$`�Libr���564@e�� �4H`ZU�SoY0t ssag�E�~� "�1�V�VLO�b/I- �pc
�`MIL;IB�mch1o Firm+�8� �b�"Acc` hXcT�PTX�;��� s Teln�0�m}B��5|��4Torqu
 imula�}�7Tou7@Pa51��Em�T_ �QC&V �ev. ocle�USB po,U � iP�a@Wd?USR EVxP+�Unexcep�tx�P�D{D{f}V�C�r�"�"�2�sV�D��j�cV�Hk u�ifoV�SP CgSUI�k��XC�6�X`Web Pl�V��9pjăa�+64.f��^ r>p�T�v�
J57À��vGrid�Qplay 76 (�X�`L&iR;�.��:K�\0ARC; 4 �120i��L#AsciiV!eRDAG�d��UplE@��� �@oCollW�Gu��� of^QޝPI  � 1�s� ��t�0tX8FK���Cy�p  2�*Porie  l�d�aFRL�1am�͉ RINT��M�I DevO0 (�&ax2 ,�0�%(}t�\rb�A/��Pa�sswo��:O"� {zes�
! �064MB DR�AM�
qG`��FR�O�� RBW��r�ciPvis�]�ByW� .�Welds ocial�4 "Pΰ�ell���mr�w�shg�s���c�XE awm��( p��v �Q��ty	 s$PR-�8�2�t!1m@-.�bo+�D�P�X��D� 2b a����r�Dr�Pb� q gged� rT1� �e8sOL��Sup��r�AR ! � OPT "W�  ���; cro�V ���SHe[�;`L�Qfq�~X�uest E��$`S��e�tex{DSp$![��P��`P@ �4YF�V�irtW�S��  ���stdpn�x�uio SWIMEST f� �F0����&�� xаߕ�51 J�����(Fr�ߕ�II)�ߓ�on��!���@M!=��RY���f>�t���mfV��լ�� �Ҍr���?���&P �3���Ҭb9����eie.T���n\@p���\R���ҭ`A���2�p����!
!�����O����7 J5����5�ӝ1Q���\ar7���XPR���k "��}���b����`P���l�nko�i���0��RAMJ����;���M������H54���js883]DER��N��Ffh�M/el���չ1d/����� �d0�/��|B�/�(  �/��<��/��p��?���.fd�/��AS9TC?��616�/��g HS|?z��as������M��?r��0�?c�r W$O��!`��%rzP]O��t\awxOV4�`�O �$�a�O�ҵ��O����O��.EN _�D�`�<_��ite_?��gv t_�� aO=%IF{?�Ԉ`���g) "s_�Epa�O�-�>n1!Ot.v$To5!�_��F���o^837�o*QogW-���o�/5-X@�PDT4B��Q�ғze�OHf4�_\7	9���MN������f�tro9?6�x�9i0���J59L��%����Ak��P����_p�o�Fp_-o0�@�?(�f1'?�pm_d��O���ٟ�O.�pe����m\�A��/_����'2.p�͆cW_��֮͠c�a/\ Ry8���(Las$����O_���0x���bo��<����e�̿"%� ���K��/?�siaf<Ϟd�?�NT+���Se����//`�C/�����'37��fiUf\����$SG���Ԁ6q��RDYaLS߱�oI�omw��_#�ps0����d�hVmj��93����E�ogW�P���ch\?�I��ퟓ� 8�o����rvi7�]�S�/������V(st�,��F���@�tl��u&5/����Td
�hWi��ݶSe��6O��sr��	��! ��y8P`��dr׏�o3PRI����a�O�/	X/��spr�ߕ��擇Li?/��3 H�6x/�d94'��6�3�q54 H�/v6353�/r4 H���&0�/�'��� X?v�72�Ie?�g13$;?��7�/58r?�'�6�/��Lo�_��t �ͅA�ϐOc�m�osK�!����O�����,�O9��O�OS�ua�lP_��8�?a_�^�g�<�_��wr+��j83�?!�_]�&��NDSO-�f7O=��!�Y�ad�O9k1l�o�s_#1�o���ip#�-Et�op�RI�N,��/I���V�A�=SE_��0�
S���Z 0+ͅcmg�Z��0 4@�"�ut[/�of��`�M�r����@�����596O_��4DЏ��U��#o(� I�c5%r_����e`���G�������c���AL"���lga33_U�oy� -<�t
��	e�@t���RTU���h�z�xo��vo;��'O�52 ����4��'�2Yu\�� vOA���42I`FĿ
d -�ݕE��� (o�[��"E3�yo��Wel�_��������WMG��Ϣ3aP@�Ϣ3wm�g[����߂�- ����On�45�?�fCqMk�IO��  �� �������1���2�g��y� R�;�Co���4(S�`�⯔��Ġ��3IF���� 1!(�z�0at��cNT��q���R8��8i5�P�82\��� O��W?��˿ݿ`￘��7��4SiZ/`<��=�K�!�cl��i5\sw/�S�AD̓��CVt�Dt.�Q�mt�_�e����V�-V�  /6��Nlo��1��\�O�/�C �/�4 �/�i`�e/�/1_��62˟2��o�/�eJ7���erv�?�) "�?�svh�?
o�N�� �?�.p[�tvshmoO�U749LO�R`r��Outl$O?�t\�?��j�_��//�/h_ mpcL��y�9\KO�j�_0�/�_�uXP�/D�cH8gO}�oOnn�O�%N�߬u�'o���np]`���oRCM�o�un�_��$./�_#��m  �H552�a�be�q38BSGR78�p�q�r0���libJ61�4�cATUP��@rmc�p545�zPsgt�r6��VCAM�3wCRI�p\rc�p�CUIF�  �q2ީptd.f�NR�EN rco�p631  - Pr�p�SCHV� Di�DOCV>aIF�L�CSUJ18�0��p1}�EIO�C  ��4�p54R�pR�`4�9�pgm�wSETf�Sta�q^�qlay,�p7�q��0MASK~�SPRXYZa�ap�7f�C�pH'OCOC��3.3�r6�p\c΂51�p���qapp.�q39�f�j50�q�us�t3�LCH��A`
?OPLG�1"��E�� "L3�MH�CR  08 (�ĀS@�Reg��C�S�p�1H��p��q5��p08\�pMDS�W  URGw�MYD���sOP��\!�MPR�ra�4�Հp!�o�f��p! p���PCM�H��R0БPath���p@aDH�ՀRm����pTP�ܠ�Հ816�50��pg��āS��ol�,�9Ղ:�FRD��p(Q�pMCN��c�c�H93�pLN=P��SNBA@�r�SHLB��֑SMnx�lrn?�63�p���q2�pL�HTC<�pX�TMILVs�r��T��PAu�Y�s�ȡTX>aEN��E-LU�th��0�@`�8�qHѰr9��`ρC95�p �Հ7���UEV��adin�(�C�����pUFRvI�eeO�VCC�p�t�VCOY���VI�P��spd�[�I�^�p�X͡tsπW�EB�p��?�HTTv�p L2�R62�p7Coo?�CG��d��IGt�
PR�I��PGSN ng��IRC��ne n��H84�prd6��R7��@�R��L�5�3�p\lcl�q8^�pD" #4�6M�� ��52�8�R6�59��|�5�r AdK�6��p��4�49��YpS��p5�̰T©qG� ML�06�pg, ��F{���ð��poJ643�pWS�pn��CLI�zdҡV��pGD����u�$�0����h�TY��<q��TO�pg���q6��-@��R5 ��OkRSY�3��68�pvģOLp�sguK�GOPIɰݠ�pS5�FR�RLP�y��S�2!�ETS1���o43 !��CP-��ryB�VRu�on�F�IPN�� Loޟ�Gene~�(S)ytE�a��I�0�����p�ytt\sg��g "�ր6q���L�yt\str�ոA�ՀA��hk_�t���yt����esؤլr��j7��moCn.�՜A��d@6���s-@�ց�yt46\�`Q���qh3��zDglli4�F�lc�`�$rt{���¥Հ��yt��w�x�U�Ӑh�8��nde��Ax�V絰����N��ͰH��epen���ytb�T��Ģ��ob3朔���h89����p���Pv�ed����4{ J7R805���0l��ձ`"t64q4����� II��d�r�p����"S��p5л%��594G��tom���!�R� J��� ��Sef3�ar3�E�t32��%�QsysG�F� ��������etr���urnk����20�x78���'��rn6�����\jftET��
jo���ta.C����gr ������� ���<���sge���017��a2�yt�yt75b����Lj(���7 �"P��T`dc ��) ��	����r�L�1%at�@O����p��daW(?�4t v/ 4oh��c8}����s?yR�?�=logm��?�;ild�?1<d �?N�@���0@O�	M���p1|O�;x@���ytV��1���O_��	8�aicC! 2�9���C��x7��6�E ��c `E?kedg?�y=wm�`ORhl$_�2G&he>�m_��M7�5l�O 24Of Oaw4OJmdh\o��;dh2���osqz�o�kl���o�oh��:��+F�et�'�-�6J8"WQ��1G (F���pDa�0��fr{F� �� ��f22.f�Fus�S�pkg�M!IN"gD�x���,��u�p�o�{��522�x�siRC�n V9M��^�992�W� ֤�J9�b�stx�'T��O 92\�6CMR/d#Z��O;��"ݎv'���tmF�����f8�vat��t�+9>e��6ft"/��z_v(��ɟ?�4o"��,���կK����vsw�8��D3ni�o��lb�� 蟮�����W�\����vsmTڴa�z�"����ο��o�f���ow�(ώ�s	lw���f���e�w�����*�vr�ys�+�N3GeN���Y25�:�oad��(Nab�NJ?��nd��� "NwV  ��@��<���rcrd�6`��le&���C�U�4;��Ok#7\��8���rk&,�F��gl��P��g�Gt��il������   P2�^���38��r� ����0���J614�A�TUPj���545�����6F�VC�AM��CRIr!7� , UIFB����2��ans��C�NRE�'��631v��RI��SCH�u�65DOCVvN�ns� CSU�T�|���0��HAE�IOC% "��5�4��R6965=\� ESET�W������7 Cuޛ MASK�t 1PRXYU�J N 7�ל�OC�O�om�513�r�,,������ ��9�8\t����]�[3�9�v!��oft�wLCH!g^�OPLG:�950ai�P]P��We f,S�r�ІCS���gW_lo��5� �p�DSW6�r70�<!Pl DKOP�P4�PRQS01� n Ad����.X#PCMAa ���0�%���vdvx; �A
TX���0��1ADIGH� �!H ,S�/r723��9AU��+ FRD!h#RM�CNr	H93��R^2SNBA"�C+ oSHLB�	SMp5�n m�J52ΑHTC���TMIL6�Se���PmO�0PA�86*�TPTX�VR�0E=LA4ool,���� P��8��\svx���qSRVT��95Q$95A\;et� UEV�@ab\AC!]�[AFR!�r��C!ol.��VCO��P��VKIP�4e�� I�t�34[SX���OWEB���@(�1T��,�l2tQ, �G�Eg\tkIGr�E#@`PPGS"��PRC�4"TANf��84��#R7��taQR�(
R5u3�tRJ68���R66a52�a- E��R65^qr Im�5a���l��573R�64q���q5`M8�RQ�CD06��,0g  �R4]0�AAWS!f9LIq%ni�@�P��SCMS�597z[M%76 J\0cTY�4L�, TO���9 (k76�f�er@R5PCO�RS�\snKR;68��CSN� ���Eq��I1Tcsn!.\0� 6��cL�EX�0[1�f��� TS1Th#@� ��P �0a �F,0VR��,QN�4{Ca
AGeneHx抳�yMG" �y<���yg_cc�y"�xcmg_�y��yGvth�yR�x3(��,�>�P�b��z1��z!� cv�yon T��yh"�xhr�x�b݉1p�`]�iA�y CV�yCP �z��x��xpt���	q�ypse��ܨ���r57� I�n���wx͉576��(p+�)� �����L� "Al��w6\�ab����j8<�B���h ��PR<�J8�zPxC;�8�J��ps��P��x96\{�(P�y�����A�xl9 � -��iv{�oR DM<�H7�z[H6�{66�3�18�x�[�tor��������y�m�!��s�Z�]�2����na�lۺ��)�޸st�K��}str��yp1sk��=�\p����^�xj932|�C��@}�)�x8R�x2}�d����.|�޸_w��.�}hk_k�FH����9!�xke*�n�9�5
���yhe�z���<,�f�l.<��H�et_w�y�"�M�c� �� �zba8k�H�Z�ent��h�\m���s����  ��d�༛�Y�;�(�PZ�@�z9Pf�yv�@ ��.������ l�n��( l�gd��=
iƋ�! Z���+�00iB\�H[�H����� -�h[�C" #���82��2�@}�O�R��� ���iB/�̿N@�"F���f���h@+�=���tk� 3OR����83�i1f�t ˚�~nc+�&�fc����5���835�z����i�;˱5:�B�ri��E�R���b݉ (ˊn�g,�@�,4�*R`ȭY�k=�mo�`�]/��p�+��ptp�z(�5\pk�=O?� ���0[ڈ��0�/�/ ? S�i�k߽�ij��0
��?�+�db���/ s50l�a��x�:��S�[d G�y�Ƌ�ce��0K�50�K1�y�6q:�Je�RDE��yqvInt�
 Pa���(�9\g{�H�91�9[�p�\:� Vi��tool<?ވ	�J[�uppK/=_��vk{��K[��Z�� Z��O�O�O�8�OK�H���?�G_rj;*h�nsdr{�H]end��Ir:�(�3��o~HC73;���/�&7;* ��{X�j�|���"�~4�  am_xOF�ve�ʘ���vI���o�?|�xj{���� �Tz{�] R5v;�J9�;989����_��p�m
�
��`����e�kR �R�}++R7�J L:;) "���Kz�/)p+zx�d	�-�|��	�633�06 �S�I~R6�st��z��:�LND��I�F K�45��-c�on{
C9�i�*a�r �jyp�	�dsc "����ENl�ey��s��l�gr��se-�
��856��`�zrpiZx=H�O4 l�^�wj��! r˛vv�:nYn�}RC:| ��� J9�Z����86-7�13J;6��8 r�JT�`�I(iR���R|"ٟc  �STD��.pLANG&�����r��ti����P���q��)0-�� E���kg
��y` ��5����R730x��(��8 (i��/ErrP��,�`���PC��x���rvg�e������8���ge@��a<����	�.���isio��ckin�� �R�(���pGi� �����؁��j	��PFK"Ƞ�XA��\@��BP�4��!��d��aa3bbPbbb������P��P��(1��SPx�Р�FS J��wJ91��685�9!	��02*4<627���Y��,����X���;s\�GFSO����sex��/�vr�����&����RG(R68'6�4����#8	G{ (� CCR���I���cc�� "�CkH���9�\�RBT}rgOPTN�4�4�2�4��?�?O"Ocrg.�8EF��8E��
8Ed޽DPN��io{n �End.�E�xa�FINT�E��7�E� n�Ea�@�E�0�"�EHQ�Ehd\mƘFHD�F��D\eCrh�F���O�Ai�E���s@BT�!Uire`�Eh�Dt�Drh�G�dCfU��ted <��-�n An�U��-�9p9�Ut2-�8-�A0E-Ęa�U�`t f �1-��2-ĥ m�U�a�U葬U-`s�U�ѬU�pB-�1�-Ā6q��U R88�U8�51_f4�`�Uticar�U�-�it� x-�l"-�MR S�f`�fTXP�U��e{pm�f" #1�fG! T�fy��fm�g���e�P�U 2�U 70�Uonjg-ĭ@._f J7�Vipp�fon,�U���X�v4.-�j79�fc��e�]h98jg�"-�\chp�WEN�vd@PNb{Sto'�� E f$�@�VgF0�el�gx��U��j8svY��f��-�6uharel�UKARo�ComTc�u�RĆL*wp\ ��V
+vY�u�fp;\e�VAN"���]k�gpcp_f1a!�I�[�f4y�wf
!� Gf Co�uairwf�FІ84_fw5 H�fH84�vo63 H�fH7�v�779_f24��7�rw69*�65�f1��g8p��V75�VI�C �f AP7v893���R0-��B�e�ck���Hs�
Ep����#fMNS+v@���VՐ�V�P_f-]��_�Q�VX�\���tcqh믅ԬU3\pSf�WT"_fdBe��Zh�in_� �03jgo�XЬU(ROB�wOG���AUe�A�^�HR�PxflRuuyQuu�g_Sf̉3uh52�3.�Ule*wriSty �6�2�6��5sv54f�4І4�0����H60�v0�h�[�08��+�=�O�a���8< ����68v�`��s�75^0��A�rw7��h�����וл�3�v3Y�7 �U �େa2f���� 29#f8�p���\ib<f���;sbs�w��o scbP1oCja��Ly2�%� -k�E"�748�V9 wf (W_�	`f��XPF���wvF�2E�X�Ϯ`we�Vp��a\wvTf͸�z;50+�"WV����B֤u��2�Y �� ���nte�g�����f04 (�gx��D��N��BPXk���I/��`o�d�@��G��apv kϥ�ib���hp
om �wfE�1A�f��Hfdn���z�8Z�f��ؿ�r�a�W�_�oi �<�al�VVAx�V�2��� 996#fVCA8��,�vast#/�q�� ��"�dp/fy�n:�fi���58�����D��odif��.e8DP��q (d��o "���o���Rg�d9Ԑ'G��st9rS���OAW���w�R73�v16"� -Rf�79�2���iTra��c�h�/�wv"TP+v̀���tpe�c�wor����+RC�59�8 S5+�809ė?��C�f�"z\�mߦ����R�E��$FL&0�p�cz�6�verv��gng_��746t�_��S_� Ch��?�� ������<th��0�89�7i3�g����%:�f!���Īx��v�� T����w&g ���rk��p��`s�H�VAGǧset99�b����$FEA�T_ADD ?	�����q�p��	x���� ��*�<�N�`�r��� ������̏ޏ���� &�8�J�\�n������� ��ȟڟ����"�4� F�X�j�|�������į ֯�����0�B�T� f�x���������ҿ� ����,�>�P�b�t� �ϘϪϼ�������� �(�:�L�^�p߂ߔ� �߸������� ��$� 6�H�Z�l�~���� ��������� �2�D� V�h�z����������� ����
.@Rd v������� *<N`r� ������// &/8/J/\/n/�/�/�/ �/�/�/�/�/?"?4?�F?X?j?|?�?�?�tD�EMO ^�y   x�=�? �?OO%OROIO[O�O O�O�O�O�O�O�O_ _!_N_E_W_�_{_�_ �_�_�_�_�_ooo JoAoSo�owo�o�o�o �o�o�oF= O|s����� ����B�9�K�x� o�������ҏɏۏ� ���>�5�G�t�k�}� ����Οşן���� :�1�C�p�g�y����� ʯ��ӯ ���	�6�-� ?�l�c�u�����ƿ�� Ͽ����2�)�;�h� _�qϋϕ��Ϲ����� ���.�%�7�d�[�m� �ߑ߾ߵ��������� *�!�3�`�W�i��� �����������&�� /�\�S�e�������� ��������"+X Oa{����� ��'TK] w������� //#/P/G/Y/s/}/ �/�/�/�/�/�/?? ?L?C?U?o?y?�?�? �?�?�?�?O	OOHO ?OQOkOuO�O�O�O�O �O�O___D_;_M_ g_q_�_�_�_�_�_�_ 
ooo@o7oIocomo �o�o�o�o�o�o�o <3E_i�� �������8� /�A�[�e�������ȏ ��я�����4�+�=� W�a�������ğ��͟ ����0�'�9�S�]� ����������ɯ��� ��,�#�5�O�Y���}� ������ſ����(� �1�K�Uς�yϋϸ� ����������$��-� G�Q�~�u߇ߴ߽߫� ������ ��)�C�M� z�q��������� ����%�?�I�v�m� ������������� !;Eri{� ����� 7Anew��� ���///3/=/ j/a/s/�/�/�/�/�/ �/???/?9?f?]? o?�?�?�?�?�?�?O �?O+O5ObOYOkO�O �O�O�O�O�O_�O_ '_1_^_U_g_�_�_�_ �_�_�_ o�_	o#o-o ZoQoco�o�o�o�o�o �o�o�o)VM _������� ���%�R�I�[��� �������Ǐ���� �!�N�E�W���{��� ����ß������ J�A�S���w������� ��������F�=� O�|�s���������� ߿���B�9�K�x� oρϮϥϷ������� ��>�5�G�t�k�}� �ߡ߳��������� :�1�C�p�g�y��� ����������	�6�-� ?�l�c�u��������� ������2);h _q������ �.%7d[m �������� */!/3/`/W/i/�/�/ �/�/�/�/�/�/&?? /?\?S?e?�?�?�?�? �?�?�?�?"OO+OXO OOaO�O�O�O�O�O�O �O�O__'_T_K_]_ �_�_�_�_�_�_�_�_ oo#oPoGoYo�o}o �o�o�o�o�o�o LCU�y�� �����	��H� ?�Q�~�u��������� ׏����D�;�M� z�q���������ӟݟ 
���@�7�I�v�m� �������ϯٯ��� �<�3�E�r�i�{���|��˽  ¸ ����)�;�M�_� qσϕϧϹ������� ��%�7�I�[�m�� �ߣߵ���������� !�3�E�W�i�{��� ������������/� A�S�e�w��������� ������+=O as������ �'9K]o �������� /#/5/G/Y/k/}/�/ �/�/�/�/�/�/?? 1?C?U?g?y?�?�?�? �?�?�?�?	OO-O?O QOcOuO�O�O�O�O�O �O�O__)_;_M___ q_�_�_�_�_�_�_�_ oo%o7oIo[omoo �o�o�o�o�o�o�o !3EWi{�� �������/� A�S�e�w��������� я�����+�=�O� a�s���������͟ߟ ���'�9�K�]�o� ��������ɯۯ��� �#�5�G�Y�k�}��� ����ſ׿����� 1�C�U�g�yϋϝϯ� ��������	��-�?� Q�c�u߇ߙ߽߫��� ������)�;�M�_� q����������� ��%�7�I�[�m�� �������������� !3EWi{�� �����/ ASew���� ���//+/=/O/ a/s/�/�/�/�/�/�/ �/??'?9?K?]?o?��?�?�?�?�9  �8�1�?�?	OO -O?OQOcOuO�O�O�O �O�O�O�O__)_;_ M___q_�_�_�_�_�_ �_�_oo%o7oIo[o moo�o�o�o�o�o�o �o!3EWi{ �������� �/�A�S�e�w����� ����я�����+� =�O�a�s��������� ͟ߟ���'�9�K� ]�o���������ɯۯ ����#�5�G�Y�k� }�������ſ׿��� ��1�C�U�g�yϋ� �ϯ���������	�� -�?�Q�c�u߇ߙ߫� ����������)�;� M�_�q������� ������%�7�I�[� m�������������� ��!3EWi{ ������� /ASew�� �����//+/ =/O/a/s/�/�/�/�/ �/�/�/??'?9?K? ]?o?�?�?�?�?�?�? �?�?O#O5OGOYOkO }O�O�O�O�O�O�O�O __1_C_U_g_y_�_ �_�_�_�_�_�_	oo -o?oQocouo�o�o�o �o�o�o�o); M_q����� ����%�7�I�[� m��������Ǐُ� ���!�3�E�W�i�{� ������ß՟���� �/�A�S�e�w����� ����ѯ�����+� =�O�a�s��������� Ϳ߿���'�9�K� ]�oρϓϥϷ����� �����#�5�G�Y�k� }ߏߡ߳��������� ��1�C�U�g�y�� �����������	�� -�?�Q�c�u������� ��������); M_q����� ��%7I[ m������ �/!/3/E/W/i/{/ �/�/�/�/�/�/�/? ?/?A?S?e?w?�?�?(�?�?�1�0�8�? �?OO1OCOUOgOyO �O�O�O�O�O�O�O	_ _-_?_Q_c_u_�_�_ �_�_�_�_�_oo)o ;oMo_oqo�o�o�o�o �o�o�o%7I [m����� ���!�3�E�W�i� {�������ÏՏ��� ��/�A�S�e�w��� ������џ����� +�=�O�a�s������� ��ͯ߯���'�9� K�]�o���������ɿ ۿ����#�5�G�Y� k�}Ϗϡϳ������� ����1�C�U�g�y� �ߝ߯���������	� �-�?�Q�c�u��� �����������)� ;�M�_�q��������� ������%7I [m����� ��!3EWi {������� ////A/S/e/w/�/ �/�/�/�/�/�/?? +?=?O?a?s?�?�?�? �?�?�?�?OO'O9O KO]OoO�O�O�O�O�O �O�O�O_#_5_G_Y_ k_}_�_�_�_�_�_�_ �_oo1oCoUogoyo �o�o�o�o�o�o�o	 -?Qcu�� �������)� ;�M�_�q��������� ˏݏ���%�7�I� [�m��������ǟٟ ����!�3�E�W�i� {�������ïկ��� ��/�A�S�e�w���𛿭���ѹ�$FE�AT_DEMOIoN  ִ����ΰ�INDE�X�����IL�ECOMP _����7����-�SETUPo2 `7�A�?�  N l�*��_AP2BCK �1a7�  �)Ҹ�ϯ�%����ΰ:�����Ե��*߹� N���[߄�ߨ�7��� ��m���&�8���\� �߀��!��E���i� �����4���X�j��� �������S���w� ��B��f��s� +�O���� >P�t��9 �]���(/�L/ �p/�//�/5/�/�/ k/ ?�/$?6?�/Z?�/ ~??�?�?C?�?g?�? O�?2O�?VOhO�?�O O�O�OQO�OuO
_�O _@_�Od_�O�_�_)_ �_M_�_�_�_o�_<o No�_roo�o%o�o�otF�z�P~� 2��*.VR�o�`* F�cLpZe�pPCx��`F'R6:��~\��{T��'��u�Q�����w�Yf*.F�
���a	�s��Ռxd�����STM ��"�-��p�Y��`�iPendant? PanelY���HO���?���[�����GIF�6�A�"�pߟ񟆯��JPG�����A���c�u�
��zJS�=��`У+���%
JavaSc�ripti���CS�Z���@���k� %�Cascadin�g Style ?Sheets�_`�
ARGNAME�.DT�lD�\@0��P�`�q��`�DISP*g�J�D�����σ����ϡ�	P�ANEL1��O�%�D�8�x�k�}�+�2 m���b���~ߐ�%�0�3��W�b�E����0�4u���b������-�(�TPEINS�.XML4���:\�H���Custo�m Toolba�r����PASSW�ORD��}nFR�S:\���� %�Password Config XoV��O��o�? ��u
�.@� d��)�M� q�/�</�`/r/ /�/%/�/�/[/�// ?�/�/J?�/n?�/g? �?3?�?W?�?�?�?"O �?FOXO�?|OO�O/O AO�OeO�O�O�O0_�O T_�Ox_�__�_=_�_ �_s_o�_,o�_�_bo �_�ooo�oKo�ooo �o:�o^p�o �#�GY�}� ��H��l������ 1�ƏU������ ��� D�ӏ�z�	���-��� ԟc������.���R� �v������;�Я_� q����*���#�`�� �������I�޿m�� ϣ�8�ǿ\������ !϶�Eϯ���{�ߟ� 4�F���j��ώߠ�/� ��S���w߉���B� ��;�x���+����� a�����,���P��� t�����9���]��� ��(��L^������� �$FI�LE_DGBCK� 1a��� ��� (� �)
SUMM?ARY.DG�hOMD:�0t �Diag Su�mmary1>

CONSLOG&�	t�CCo�nsole lo�g�=	TPACCN�/%�4/?�TP Acco�untin�>
�FR6:IPKD?MP.ZIPh/l�
�/�/@P Exc?eption�/n+�MEMCHEC�K*/�@?�M�emory Da�taA?�LN�)	FTP��?'?��?K7�mmen�t TBD�?u7 �>)ETHERNET�?f�!O�HOCEther�net �fig�ura�/D�1DCSVRF�?�?�?�O�Q1%�@ ve�rify all��O�M,��EDIFF�O�O�OO_R0�%�Hdiff�Q_W�!�@CHGD�1F_-_?_�_ Xf_�_S+P�Y2�_8�_�_Xo �_ooGD3No5oGo�o� no�fUPDATES."p�iFRS:\� a}DUpda�tes List�afPSRBWLOD.CM�hLr��c�PS_RO�BOWEL�?<>�aHADOW�o�o��of�Q3Shad�ow Chang�esi��=�&�NOTI�OA�S���O5Notif�icqB���O�AJ?�nc��p��� D��L��󟂟��� ;�M�ܟq� �����6� ˯Z��~���%���I� دm�����2�ǿٿ h�����!�3�¿W�� {�
ψϱ�@���d��� ߚ�/߾�S�e��ω� ߭߿�N���r��� �=���a��߅��&� ��J���������9� K���o����"����� X���|�#��G�� k}�0��f ���,U�y ��>�b�	/ �-/�Q/c/��// �/:/�/�/p/?�/)? ;?�/_?�/�?�?$?�? H?�?�?~?O�?7O�? DOmO�?�O O�O�OVO �OzO_!_�OE_�Oi_�{_�$FILE_�LpPR[p���_P�����XMDONLY �1a�UZP 
 �
_�_._oR_o ;o__o�_�o�o$o�o Ho�o�o~o�o7I �om�o� ��V �z�!��E��i� {�
���.�ÏՏd��� �����*�S��w�� ����<�џ`������ +���O�a�🅯����8���߯�ZVISB�CK�X�Q�S*.�VD�0���FR�:\��ION\DOATA\�â���Vision VD file\� j�����̯ڿį���� �4�ÿX��|ώ�� ��A���e�w�ߛ�0� B���f��ϊ�ߛ��� O���s����>��� b�����'����� ������'�L���p� �����5���Y���}����$�ZMR2_G�RP 1b�[�C4  B� �	 �Qk}h E��� E�  F@ F�5U��/
h L���M���Jk�K��v�H�,�Hk{��?�  ��/h 9tQv8���6h�%��A�  3EBMHeB�a `�E	@i/g��h /@UUU�U���>�]�>П���;r8	=�==E��<D��><�ɳ<�����:�b�:/�'79�W�9
�@�8�8�9��T/�Q/�/e�E7� E?p �D�D�/�D�  D�  Cζ/�9
_CFG c�[T �/?0?|B?�NO �Z/
F0x1 }0��RM_CHKTY/P  �P� �P��P�P��1OM�0_�MIN�0
����0�PX�PSSB��#d�U�P�i�?	�3O$O�UT�P_DEF_OW�P
�Y?AIRC�OM�0JO�$GE�NOVRD_DOr�6�RxLTHR�6� d�Ed}D_EN�BiO }@RAV�CGe�7� ���FnH E��� Ga H��� H�@Jh!`�/O?_�G_X_n{ ��AOU�@-kN {NB{8���_y_x�_�_�_  C�� �	$o�XYoilCOmB���AVb~	�Y+O�@SMT�Cl�IZ �04d�$HOSTC�"{1m��k 	
x
{
2:byeV� ����zu� ���$�GH��p	ano?nymousK�y� ��������	- �A�c�V�h�z��� ���ԟ����M� _�@�R�d�v���ˏݏ ����7��*�<� N�`�����������̿ �!�3��&�8�J�\� ����ïկ׿����� ���"�4�w�X�j�|� �ߠ����������� �0�sυϗϩϫߜ� �����������K�,� >�P�b���s��ߪ��� ������G�Y�k�L �p������ � $6YZ�� ~����	�- ? /SuB/h/z/�/ �/��/�/�/�/
?-/ _qR?d?v?�?�?� �//?�?I/*O<O NO`OrO�/�O�O�O�O �OO3?E?&_8_J_\_�n_�g�aENT 1�n�i�  P!\�O�_  �@�_ �_�_o�_+o�_Ooo [o6o�o�olo�o�o�o �o�o9�oo2 �V�z���� �5��Y��}�@�v� ����׏�������� +��T�y�<���`��� ��埨�	�̟ޟ?���c�&���J�QUI�CC0��p�!1�72.8.9.225����1���ү�3���24������!ROUTER���`�r�ӿ!PCJ�OGԿ��!1�92.168.0�.10����CAMgPRT$� �!�11�K�2�RT��O��a��ψTNAME �!�Z!ROB�O=���S_CFG� 1m�Y ��Auto-started�4/FTP�?[��? �O��O�߼������� �O�(�:�L�o�]������������#� �:4�F�X�9�l��P� ��������z������� #F���Yk}�p���?�=SM�65233)�
= _�,Rdv�K�`����  %���5/G/Y/k/}/""q��?�?�?�/3 ?&?8?J?\?/�?�? �?�?�?�/m?�?O"O 4OFOXO�/�/�/�/�? �O?�O�O__0_�? T_f_x_�_�_�OA_�_ �_�_oo,ooO�O�O Eo�_�o�O�o�o�o�o �o(:L^�o� ����� �Co UogoH�{�o����� ��Ə����� �2� U�׏U�z������� ��)�;��O�q�R� d�v�����]���Я� ���)���<�N�`�r��������_ERR �o�ʡ���PDU�SIZ  3�^�L��ȴ>�WR�D ?"��� � guest-�!�3�E�W�i��{���SCDMNG�RP 2p"�˰��3���-�K�� 	P0�1.05 8�� ������> j W 2�1�� ꛿ ���T�����������/����$���Ͽ�Q�<�u�`�������  � � 
��N(�P�,�(����Q�����������l�� 8�#{�d������"ߙ�_GR�OU��q����ҍ�	����4S�QU�PD  �ȵ�X��TY������TTP_AUT�H 1r�� <�!iPenda�n����8�g�!�KAREL:*8����KC-�=��O�%�VISION SETb�����!������"� �� _6H�l~���CTRL s������3���F�FF9E3���FRS:DEFA�ULTFA�NUC Web ?Server�� ��	�Ĵ}��������WR_CONFIG t��� ��IDL_CPU_PC*�3�B��I  BH/%MIN:,��M%?GNR_IO������Ƿ1 NPT_S_IM_DO&�+�STAL_SCR�N& ��*TPM?ODNTOL�'�+bRTY�(I!�&��N��ENB�'��-$OLNK 1u���Q?c?u?�?�?�?|�?52MASTE~ ���52SLAVE �v��34��O_C3FG�?IUO��O>BCYCLE>OD�$_ASG 1w����
 �?�O�O �O�O�O�O__1_C_�U_g_y_�_�;tBNU�M�Ĺ
BIP�CH[O��@RTRY_CN*�"ĺBP�!���P1�ȵ B;@Bx�>�Jo��1 SDT_ISO�LC  ��f��$J23_DS4��:��`OBPRsOC?�%JOG^��1y�;��d8�?��[�o�_?؟֟O|QNs���V����-��~o�h�`Y A�_�bP�OSRE�o�&KANJI_�0���/k�~+�MON zg��2�y�Ϗ�����Ҿ)�0c{,�09�T���e�_LY �R��_k�EYLOGG+IN@����ȵ��$LANGU�AGE k2e$ 㑱�LG1bY|�2���3�x��ʗ���O � '�0,�� �
q��3�MC:\�RSCH\00\���LN_DISOP }�?f�M�Km�OC�"@"Dz�h#�A�OGBOOK ~K��w�0��w�w���X��� -�?�Q�c�u���11����	���h��޿����ॐ_BU�FF 1@= ���)�����E� a�sϠϗϩ������� ���B�9�K�]�o���ߓߥ��ߜ��DC�S �� =��͗�ֿM�l:�L��^�p���IO 1��K No����� �����������%� 9�I�[�m��������� ��������!3E�Y��Ex TMlnd ������ 0BTfx��� ����//����SEV`}��TYPln��/�/�/)-P�RS�P���b�FL 1���`��?,?>?P?b?t?��?�/TP��loq">��NGNAM�d���Ւ��UPSu�GI��U\�e�1_LO{AD�`G %}��%DF_MOT�N$�FOݠMAXUALRM�Wk�X\@N�1_PR�T`ԣ4��Z@Cx��ꩦ���OV�9ŜC�`P 2]��K �9�	q!�P]  � �OQ�R9_$_6_o_� ]_�_�_�_�_�_�_�_ oo@oRo5ovoao�o }o�o�o�o�o�o* N9rUg�� �����&��J� -�?���k�����ȏڏ �����"���X�C� |�g�������֟���� ݟ�0��T�?�x��� m�����ү��ǯ�� ,��P�b�E���q����SGD_LDXDI�SA�0�;��MEM�O_AP�0E ?=�;
 j �� ��*�<�N�`�rτ�~Z@ISC 1��; �����T�A����ϛ�$��Hߙ�C_MSTR �B-~g�SCD 1����<߶�8��������� "���X�C�|�g�� ������������	� B�-�f�Q���u����� ��������,< bM�q���� ���(L7p [������ /�6/!/Z/E/W/�/ {/�/�/�/�/�/�/? 2??V?A?z?e?�?�?��?X�MKCFG ��vݽO�CLTAWRM_�2��G�B� P�2�@>OFD{@M�ETPU�C�@���~�ND�@ADCO�L`E�@kNCMNT�O tEo� ��v��N5C.A�O�DtEP�OSCF�G�NPgRPM�OYST@{1��� 4@��<#�
oQ�1oU_ �Wk_�_�_�_�_�_�_ o�_oOo1oCo�ogo�yo�o�o�o�o�atAS�ING_CHK � �O$MODA�QC��?���>+uD�EV 	��	�MC:_|HSIZ�Eѽ���+uTAS�K %��%$1�23456789� ��u)wTRIGW 1���l#E%�̀)����S�6�%C�vY�P�q>�At*sEM_INF 1�#G� `)�AT&FV0E�0`�׍)��E0�V1&A3&B1�&D2&S0&C�1S0=ƍ)A#TZ׏+��H/�W��K���A����j�ӟ����	� ��.�� �����;����Я ⯕����*�<�#�`� �%���I�[�m�޿� ���K�8����n�)� ��y϶���{��ϟ��� ÿտF���jߡ�{ߠ� S������������� ��T���+ߜ��a� ��	�����,���P� 7�t���9��]�o�� ����(:q�^���=����XN�ITOR�@G ?�s{   	EOXEC1�32%3%4%5%�p'U7%8%9�3  ��$�0�<� H�T�`�l�Px���2�2�U2�2�2�2�U2�2�2�2��3�3�30+qR�_GRP_SV �1��� (�a>������*��=E�����4�X>��Z}ƶq_D{�~�1PL�_NAME !�#E0�!De�fault Pe�rsonalit�y (from �FD) �4RR2��! 1�L68�L@�1P
d d�?v?�?�?�?�? �?�?�?OO*O<ONO `OrO�O�O�O�O�O�OJx2e?_ _2_D_V_@h_z_�_�_�_r<�O �_�_�_o"o4oFoXo@jo|o�o�o�i�V�_"�n
�o�oNtP�o* <N`r���� �����&�8� n���������ȏڏ ����"�4�F�X�j� |�K�]���ğ֟��� ��0�B�T�f�x���𜯮���Ү F�nH F�� G�=��'�   �����"d���0�B� &�d�r��׭Ҫ\���p����ݿ� ͸ ��� ��0�6�T�v�� �ϩ�ͰA�  ��˿��Ǹ]0�� �ƿ3�¿W�B�{ߍߐx߱�B5K3�9^0�`�!0 � ��0�� @D��  ��?����?x� ��!A����x�$��(;�	l��	 ���p�V� ]0M� � � � �l���r� K(��K�(�K ��J��n�J�^J&Ǔ�2�������� @Y�,@C�z@I�@��������N��o��f���_�I���SѬ�Ä��  <��~% �3�������!?s8y�
�}/�!�x����T� ܌��������}��  �  ������7  ����������	'� �� 0I� ��  �����:��ÈTÈ=��1�l��	�(|�� ���Ѧ���ψ��N@0�  '����@2��@Ϙ��@!����@�)��C@0C���\CI�CM�CQ��� ��� .� O %�~���� ���B���@0��l@� ��!Dz���V��//+/Q/���� �H@q)q�%�  ����  �� p�!?�ff0���/�/V/ ���/;��8� !?/:��D4�� \6Pf8�)c�\�\��?Lv �$���;�Cd;�pf�<߈<��.<p��<�?L:D��ݧA���d��|��?fff?��?&@��@��� B�N�@T� ,E�	��	A���dO �O�7H��/�O�O�O �O _�O$__H_Z_E_~_�MEF�m_�_ i_�_UO�_yI�_2o�X�C��E��"Gd G;ML!o�omo �o�o�o�o�o�o�o$ H��iww9��_ �o�U��*�<�ڪ����/�6�������ď��菎�A�A�����C؏=�ԏ��X��񨑟,���>��  �P��"@�z<��E� C���s��x�؄�(������/�B�/B"��}A��#A���9@�dZ?v�ȴ,��~���<)�+� =��G��j���q����
AC
=�C��������� ��p�C�c�¥�B�=���ff��{,�I����HD-�H�d@�I�^�F8$ �D;ޓܪ�̠J�j��I�G?�FP<����QpJnPH��?�I�q�F.� D��Ɵg�R� ��v��������п	� ��-��Q�<�Nχ�r� �ϖ��Ϻ������)� �M�8�q�\ߕ߀߹� �߶��������7�"� [�F�k��|����� ������!���W�B� {�f������������� ��A,eP� t������ +;aL�p�����(����3�:��1��%�3��V��/"��(/:/�!4M��xT/f/F1�=Ӏ/��/4Ue'��T9�-�)�/�/?�/4?�"<]�P�2Pf>�q ��?��?�?�?�?�9���(�?�?/OO0?OeOPO�QB�hOzO �O�O�O�O�O�?t.__R_@[/X_b_�_`�_�_�_�_�Q{f�_��_o
o@o.odorj  2 FnH"��F��"�G=��B# ��C9)��@|��@��o �q�o{E��� F��`�H C�����oA`�m�kE�0wGa�O����{?ސ�q ��\d  zq: `�
 �!� 3�E�W�i�{��������ÏՏ�������q ���P+�~Y���$MSKCFMA�P  �%� ^f�q�qp��D�ONREL  �X5[��0D�E�XCFENB��
8Y����FNC�����JOGOVLIMҍ�d����dD�KE�Y�����_P�AN����D�RU�N��SFSP�DTYw0������S�IGN����T1M�OT럜�D�_C�E_GRP 1��%[�\�O��O �&��d�Q��u�,� j���b�Ͽ��Ŀϼ� )�;��_�σϕ�L� ��pϲ��Ϧ��%�� I� �m��fߣ�OvD�QZ_EDIT���U��TCOM_C_FG 1�Q������"�
��_AR�C_��X5ؙT_MN_MODE���縙UAP_C�PLF４NOCH�ECK ?Q� W5�H������ ����'�9�K�]�o������������v�NO_WAIT_L��l�׾�NT���Q�z�{_ERRȡs2�Q��1� ��t���H*���Ԛ�`�OI�Px �
F��A6y��犑������u��=/��@���I8�?0|4��pdB_PARAMJ�Q����߷�7so�� =�`345678901�/ * �?/Q/-/]/�/�/u/0�/�/�+�7�?<��7?��UM_RSPACEN��$�p?�z4�$ODRDS�PE㌦��OFFS?ET_CAR�Ќ�έ6DIS�?�2PE?N_FILE�0��$��֌1PTION�_IO
��@M_�PRG %\:%�$*IO[N�3WOR�K �Χ�� ����FQtҡ�r�^�(�d�@(7�A	� ��x�A5��c���0RG_DSBL'  \5���|_��1RIENTTO��9�C��pZ��a��0UT_SIM_EDGX�+��0V�0?LCT �%��x�Dx=gT_PEXh���?�TRATh� d��T�0UP )�u^�Ӡ�ooX�_:oHi�$�2ǣ��L68L@}�_S
d d'? �o�o�o�o�o�o�o 1CUgy��@�����I2~o '�9�K�]�o���������ɏ9�<���� )�;�M�_�q������� ��H�j3�H1`��XRP�C�U�g�y� ��������ӯ���	� �-�?�Q� �2����� ����Ͽ����)� ;�M�_�qσϕ�d�v� ��������%�7�I� [�m�ߑߣߵ�����X�ϡ��*��S�H�Z�?�}����@��&?������� �����+�I�O�m�����?@�����A�  ������� ���M8q\�����z�d`O�P1��k����sd`�B0 ���D$@ @D�C  DD?Q�D	��E� � ;�	l1	 ���p�s& ' j � _� � ʉ��� H<zH<W��H3k7G��CG���G9|�+c	�H
��� CC9P/9P49S;Q9�/��9  ���  1!�H7 3�����/1/C/�BY����XQ��^�H�<Pq/ ܩ/�"2�#�3�.��    ��0�� �  0�6�/?�	'� � M2�I� �  ����
=���q?�;�&��@&�/ ��A�?4;�B�?r�NEPO  'VP�3D�b CEPC��+\Cf Cj Cn/@O|ROߑ  ���~�D%%���� �B`���FEP�E˜@XP�E5z�_s/8_#_�H_n_��� ��H]2�Y�A�U  ��C�H�A�0p�Q?�ff���_�_�s_ ��o(k�18 �0>oLj-�!adTW�0yfP�h�Y�yy�3�?L�0�T�;�C�d;�pf<���<��.<p���<�?ij��WA��Eل1d�31��?offf?�@?&+p�VT@��=r�N�@T�IuՉ�� &q-�0!��w e o������ A�,�e�w�b������� я����l���O���CE���2Gd G;�|>��� ��ß���ҟ���� A�,�e�����V��� �د6���r�#�5�G�Y��Z� �_�f���@����̿��A @!A�@%���5�C��Z�x��/i�?�؈�p���ϳ�U�P��2�]!YNE� CU%�̣�Ŀ����E��@I�!t�B�/�B"�}A���#A��9@�d�Z?vȖ+~��~���<)�+?� =�G�(߇����q���
A�C
=C������녡� ���p�Cc�¥��B=��ؿff�{��I����HD-�H��d@I�^�F�8$ D;���ڭ�̠Jj��I��G�FP�<��QpJn�PH�?�I�q�F.� D��E �τ�o�������� ���&��J�5�n�Y� k������������� �� F1jU�y ������0 T?xc��� ����//>/)/ ;/t/_/�/�/�/�/�/ �/�/??:?%?^?I? �?m?�?�?�?�?�? O �?$OOHO3OXO~OiO@�O�O�O�O�O��(}�ϳ�3:�O�a��<)U�E3�V�_+_�9R�E_W_t�4�M��q_�_t��=�ӝ_�_4Ue'��T9�]�Y	o�_�-ooQo?lz�P�bP�n�����o�O�o�ox�o�i���(�L7\�mt�B����������o��K�9�o�]�/ u������ŏ�ُ�{f��9�'�]�K������  2 F�nH��F�Щ�G�=��B@P!�.�C9F��p��@2���	��~C�E�� F����H C���S�b����������¯Dԯ��?����y��C�C�|�C�}�
 ۯ>�P�b� t���������ο�����(ϧ�� ���m[�~Y��$P�ARAM_MEN�U ?�U��  �DEFPULSE�4�	WAITT�MOUT��RC�V�� SHE�LL_WRK.$�CUR_STYLv����OPT�N��PTB����C��R_DECSN�� teG�A�S�eߎ߉ߛ� ������������+��=�f�a�SSREL?_ID  �U�a��u�USE_PR_OG %p�%b���v�CCR����a�x���_HOST !p�!�����AT�`��8����:�|t���_TIME������a�GDEB�UG��p�v�GINP_FLMSK�����TR����PGA��� ��{�CH�����TYPEm�y�a�[���� ��!JEW i������� �"////A/j/e/w/ �/�/�/�/�/�/�/?�?B?��WORD �?	p�
 	�RS��	�PNS2u��~2JO�
��TE[��?CO�Lu>8�?>L�� ��P��p���TR�ACECTL 1��Uz� .��{ ������|1LFDT Q��U�^@#@D � �sc01A kH�s@��BP��B��B�D�DU	�D
�D�s@��{O�O�O�O�O �O�O�O__/_A_S_ e_w_�_�_�_�_�_�_ �_oo+o=oOoaoso@�o�o�o�o�j�a�d �o $6HZl ~������q/ kEC�U�g�y��� ������ӏ���	�� -�?�Q�c�u������� ��ϟ����)�;� M�_�q�����gI���� ӯ���	��-�?�Q� c�u���������Ͽ� ���)�;�M�_�q� �ϕϧϹ�������� �%�7�I�[�m�ߑ� �ߵ����������!� 3�E�W�i�{���� ����������/�A� S�e�w����������� ����+=Oa s�������� '9K]o� �������/ #/5/G/Y/k/}/�/�/ �/�/�/�/�/??1? C?U?g?y?�?�?�?�? �?�?�?	OO-O?OQO cOuO�O�O�O�O�O�O �O__)_;_M___q_ �_�_�_�_�_�_�_o o%o7oIo[omoo�o �o�o�o�o�o�o� EWi{��� ������/�A� S�e�w���������я �����+�=�O�a� s���������͟ߟ� ��'�9�K�]�o��� ������ɯۯ���� #�5�G�Y�k�}����� ��ſ׿�����1� C�U�g�yϋϝϯ��� ������	��-�?�Q��c��$PGTRA�CELEN  �b�  ���a��w�_UP �����љ�В���w�_�CFG ������a������������׉���DEFSPD ����`щ��w�IN~��TRL ������8�F�PE_C�ONFI�Ш��O������WLID�ө��	��LLB 1���� t�?B�  B4��� ��� ����� 88�?�0�K�0�G�i�k�}� ������������5Ak��� ��2��	�?~��GRP 1����lb�A�  ��333a�A���D�@ D�� �D@ A@�Ta�d+������� 	='����#´#��B 9!�///O/9/s/
?��?����/�/��.�/ =o=	7L�/?�/?P? ;?t?_?�/�?�??�?<�?�?  DzC Oa�
OHO�?XO~OiO �O�O�O�O�O�O_�O�_D_/_h_S_�_�Z!�a�
V7.10�beta1�� �Ax���R�y�y�Q?���Qo>�\)�QB0����PA��SBp���QA�9Sy�b
a�S �_2oDoVoho��Ap���"���o��o�o�o�Ҹө�KNOW_M  �|�֦�SV ���/���5O8 J\u_�k}��Ҕ���M]�z�Д��R	��%%��"��|���G� ��u��P@��a�]�a�q�m��`��MR]��}��&%O�P��$ӏ�KST]1� 1���
 4 ��vi�Q:��"�4�F� w�j�|�������ğ	� ���?��0�u�T�f� ���������ү���2� �a��<K��^35�G�Y�k���4���������5 ۿ�����6.�@�R�d��7�ϓϥϷς�8������
��M_AD  �����OVLD  ���G�PAR?NUM  ���߾��T_SCHy� ���
�����0�U�PD��������_CMP_�p|�pp�'�e��ER_C;HK�����j�⌝��RS��oW_#MO{���_��տ_RES_G�� � o����������� ����2%VI@zm`�R�4�\�l� �Q������S�ڰ �S�-�9X] S��x��S���� ��S�&��//S�V 1���a�q�@c?\�THR_INR��~��r�e�d�&MASS�/ �Z�'MN�/�#MO�N_QUEUE C���f"��a��N��U��N�&��0�END1;�79EX1EF?75\�BEE0'?>3OPTIO$7D��0PROGRAM7 %�*%0T/���2TASK_I�{ԍ>OCFG ��/���?"@DAT5A�s�+K��"�2��O�O�O�O�O�O �O_!_3_E_�Oi_{_x�_�_ROINFO�s�oM�
4[_�_
oo .o@oRodovo�o�o�o �o�o�o�o*<�N`�W�T�oL ؊	!A�K_%A�8+I�^�vENB|б}�)��v2��xG%A2���{ P(O8�4�F� C�e���z_EDIT �+O����DWER�FLg8|# �RGA�DJ ��:A����?"���!߆1��q�]��3?���A<@��v�%<�l�ӈ���q2Y�)��R	H0le��{"6�?
��A�F$�t$ܖ*z�/� **:�� "�����d�1�f�Ցd�[�_"U�#���3� E�s�i�{�������߯ կ�a���K�A�S� Ϳw���������9�� ��#��+ϥ�O�aϏ� �ϗ�߻�������� }�'�9�g�]�o��ߓ� ��������U����?� 5�G���k�}���� -����������C� U���y��������� ����q-[Qc ������I� 3);�_q���t&	>O@/Հ./ g/R$ݙ�/ߓU/�/Q/��/�/�PREF S�)�ՀՀ
߅?IORITY�72F}��MPDSP�1�яG7UTFǓކOoDUCT
A�:��/��OG��_T�G΀B���2TOE�NT 1� �(!AF_IN�Eq0OG!t�cpO6M!u�d%O^N!ic�mMOu��2XY"��v���X1)� ��O�OX0��O�O�E �O)__M_4_F_�_j_ �_�_�_�_�_o�_%o7o*�3"��=Y�yo��o��>��J�B�/�io�o��������AK�,  �0�q'9K]X5��7�pHANCE C�)��rrn{d�o��uyw	3�?"3ق��PORT_NUUMr3X0����_CARTREP�R0����SKSTAvq7 C�LGS @�ȍ��K�X0U�nothing �����̏܌������#��?k�TEMP �ɕ94����_�a_seiban �/���/��͟���ܟ � �9�$�]�H�Z��� ~�����ۯƯ���� 5� �Y�D�}�h����� ſ��¿����
�C� .�g�R�wϝψ��Ϭ� ����	���-��*�c� N߇�r߫ߖ��ߺ��� ���)��M�8�q�\����6�k�VERSI�P0�7�� d?isable�r<�SAVE ʕ:�	2600H8K44����,�!�0.�@�_Od� 	��{2$ /����X�e����	-;
��c�n� ��L��_�0 1˧K�� "����0URGEpB�0T6>5�WFF� DOr6�r�6W�0��"�WRUP_�DELAY ��;�R_HOT �%%&~1��+R_NORMALy�2���SEMI��"/�!QSKI%P���w�x��g/ ��/�/�/r-�5�/�' �/??(?�/L?:?\? �?�?�?l?�?�?�? O O�?"OHO6OlO~O�O VO�O�O�O�O�O_�O 2_ _V_h_z_@_�_�_��_�_�_�_���$R�BTIF?�RC_VTMOUT�B���`DCR�ϾE) �~!A����DA��D�+�w�b�F7��r-������,���_���~A˷����r/�o�/ ;�C�d;�pf<���<��.>�]�>П��o��o'8} 8^p ������� ���$�1%RDIO_TYPE  ��.�EFPOS1� 1���  x�����Ώ��� {����:�Տ7�p�� ��/���S�ܟ��� ՟6�!�Z���~���� =���دs����� ��� D�V���=�����¿ ]�濁�
ϥ��@�ۿ d�����#ϬϾ�Y�k� �����*���N���r� �oߨ�C���g��ߋ� �&������n�Y�� -��Q���u������ 4���X���|���)�;� u�����������B ��?x�7�[ �����>)b ��!�E��{ /�(/�L/^/�/ E/�/�/�/e/�/�/? �/?H?�/l??�?+? �?�?a?s?�?O�?2O �?VO�?zOOwO�OKO �OoO�O�O_._�O�O _v_a_�_5_�_Y_�_ }_�_o�_<o�_`o�_x�o�o|�2 1ш� 2oDo~o�o�o &oD �ohe�9�] ��
�����d� O���#���G�Џk�͏ ���*�ŏN��r�� �1�k�̟��🋟� ��8�ӟ5�n�	���-� ��Q�گu�����ӯ4� �X��|����;��� ֿq�����Ϲ�B�ݿ ��;Ϝχ���[��� �ߣ��>���b��� ��!ߪ�E�W�iߣ�� ��(���L���p��m� ��A���e������� �����l�W���+��� O���s�����2�� V��z'9s� ����@�= v�5�Y�} ���</'/`/��/ /�/C/�/�/y/?�/ &?�/J?�/�/	?C?�? �?�?c?�?�?O�?O FO�?jOO�O)O�O�o�d3 1ҵo_OqO �O)__M_SOq__�_ 0_�_�_f_�_�_o�_ 7o�_�_�_0o�o|o�o Po�oto�o�o�o3�o W�o{�:L^ �����A��e�  �b���6���Z��~� �����Ə �a�L���  ���D�͟h�ʟ��� '�K��o�
��.� h�ɯ�������5� Я2�k����*���N� ׿r�����п1��U� �y�ϝ�8Ϛ���n� �ϒ�߶�?������� 8ߙ߄߽�X���|�� ���;���_��߃�� ��B�T�f�����%� ��I���m��j���>� ��b����������� iT�(�L� p��/�S� w$6p��� �/�=/�:/s//��/2/�/V/�/�O�D4 1��O�/�/�/V? A?z?�/�?9?�?]?�? �?�?O�?@O�?dO�? O#O]O�O�O�O}O_ �O*_�O'_`_�O�__ �_C_�_g_y_�_�_&o oJo�_no	o�o-o�o �oco�o�o�o4�o �o�o-�y�M� q���0��T�� x����7�I�[����� ����>�ُb���_� ��3���W���{���� ��ß��^�I������ A�ʯe�ǯ ���$��� H��l���+�e�ƿ ��꿅�ϩ�2�Ϳ/� h�ό�'ϰ�K���o� �ϓ���.��R���v� ߚ�5ߗ���k��ߏ� ��<�������5�� ���U���y������ 8���\�������?� Q�c�������"��F ��jg�;�_����/45 1�?���n� ��f���%/� I/�m//�/,/>/P/ �/�/�/?�/3?�/W? �/T?�?(?�?L?�?p? �?�?�?�?�?SO>OwO O�O6O�OZO�O�O�O _�O=_�Oa_�O_ _ Z_�_�_�_z_o�_'o �_$o]o�_�oo�o@o �odovo�o�o#G �ok�*��` ����1���� *���v���J�ӏn��� ���-�ȏQ��u�� ��4�F�X����ޟ� ��;�֟_���\���0� ��T�ݯx�������� ��[�F�����>�ǿ b�Ŀ����!ϼ�E�� i���(�b��Ϯ��� ��ߦ�/���,�e� � ��$߭�H���l�~ߐ� ��+��O���s��� 2����h�������x9�16 1�< ����2����������� ����R��v �5�Yk}� <�`��� �U�y/�&/� ��/�/k/�/?/�/ c/�/�/�/"?�/F?�/ j??�?)?;?M?�?�? �?O�?0O�?TO�?QO �O%O�OIO�OmO�O�O �O�O�OP_;_t__�_ 3_�_W_�_�_�_o�_ :o�_^o�_ooWo�o �o�owo �o$�o! Z�o~�=�a s�� ��D��h� ���'���]�揁� 
���.�ɏۏ�'��� s���G�Пk������ *�şN��r����1� C�U����ۯ���8� ӯ\���Y���-���Q� ڿu�����������X� C�|�Ϡ�;���_��� �ϕ�߹�B���f�L�^�7 1�i��%� _�������%���I� ��F����>���b� �������E�0�i� ���(���L������� ��/��S��  L���l�� �O�s�2 �Vhz�/ /9/ �]/��//~/�/R/ �/v/�/�/#?�/�/�/ ?}?h?�?<?�?`?�? �?�?O�?CO�?gOO �O&O8OJO�O�O�O	_ �O-_�OQ_�ON_�_"_ �_F_�_j_�_�_�_�_ �_Mo8oqoo�o0o�o To�o�o�o�o7�o [�oT��� t��!���W�� {����:�Ï^�p��� ����A�܏e� ��� $�����Z��~���� +�Ɵ؟�$���p��� D�ͯh�񯌯�'�¯�K��o�
���yߋ�8 1ז�@�R���
� ��.�4�R��v��s� ��G���k��Ϗ�߳� �����r�]ߖ�1ߺ� U���y�����8��� \��߀��-�?�y��� �����"���F���C� |����;���_����� ������B-f� %�I��� ,�P��I� ��i��/�/ L/�p//�///�/S/ e/w/�/?�/6?�/Z? �/~??{?�?O?�?s? �?�? O�?�?�?OzO eO�O9O�O]O�O�O�O _�O@_�Od_�O�_#_ 5_G_�_�_�_o�_*o �_No�_Ko�oo�oCo �ogo�o�o�o�o�oJ 5n	�-�Q� ����4��X�� ��Q�����֏q��� ������T��x�����7�������MAS�K 1�û������XNO  ����MOTE�  3����i�_C�FG �p������PL_RANG�l�g�t�POWER� �õݠ|�S�M_DRYPRG %p�%m���TART �ծ�#�UME_PRO������_EXE�C_ENB  zd�x�GSPDX�우����TDB̽�ϺRM޿ϸI_�AIRPUR�� �p�B�<�ٛMT_��TРn��OB�OT_ISOLCB1��8�����9�z�NAME p��n�ۙOB_OR�D_NUM ?�ը5�H8�44 g���bҘ ����/(/�^/�Ҧ/���P�C_TIMEOU�T�� x�S23�2��1�4�γ �LTEACH PENDANP�X��������l��j�Mainte�nance CoKnsg��߾�"���f�No Use ���߮���0�B�T��h�NPO2�RҤ��z�e�CH�_L[��p���	����!UD1�:���R�VAIQL��R����x�e��PACE1 2�p�
 �濫��{鋓������9˺�?8�?�%��� %���4IDu� ������Y����� �):!4�8�Uu ������/ �):/!/O/q�� �U/���/ ?�/? 6??K?m//�/�/�/ c?�/�/�/�?O2O	O Oi?{?�?�?�?_O�? �?�OGO_._@_'_eO wO�O�O�O[_�O�O�_ o�_+_<o#oQos_�_ �_�_Wo�_�_�o�o 8Moo�o�o�o �o�o�o�D��4� �I�k}���a� ��돽��0�B��+�X�2a�s����� ��W�͏�����4�U�<�j�o�3~����� ��Ɵt����<��� Q�r�Y���o�4���� ��ѯ㯑��)�8�Y�@�nϏ�vϤ�o�5�� ʿܿ� Ϯ�$�F�U߀v�9ߋ߬ߓ���o�6 ����������A�c� r��V�������o�7����(�:���^� �����s���������o�8�!�3�E�W� {���������o�G �/� m�
u d  /��� ���/Nl -S -L/�/p�d� z ��/�/�/�/??&? /./@.1:n?�;�?�/ �/(?�?�?OO*O<O 2?D?V?h?�?�O�O�? �?HO__&_8_J_\_�ROdOvO�O�O�_ ` @p��U]/ o�O�IAakU�_Ro doj_DjEowo�o�o�o �o�o%�o�o= ASe���	� ��3�E���+�]����a�o\
#o�o�_MODE  /^
�S �/��_�Z�oH������	��㟐�CWOR�K_AD�
�O�4��R  /�< 1���_INT�VAL�a�%�R_OPTIONR�� %���V_D�ATA_GRP �2�uX:D�@P П��̟�˩͏��� 1��U�C�y�g����� ��ӿ������	�?� -�O�u�cϙχϽϫ� ���������;�)�_� M߃�qߧߕ߷����� ���%��I�7�Y�[� m����������� ���E�3�i�W���{� ������������/ SAwe�����P�$SAF_DO_PULS��Q�A��� CAN�_TIM��E}��R ���Ƙ�qsy�֡��Yo�K�C կ����� �l//%/7/I/[/Ve��C�2�$$K�)d�$�!ѢIf)�P5��/�/�/���)�/ ��4�w_ �R  T0��!?^?p?�?�9T D���?�?�?�?�?  OO$O6OHOZOlO~O �O�O�O�O�OU�s��'�O$_6_�I�  �T;��o��WQo�p�M
�?t��Di��[~=Z0 � �� o�[Q[SC�_�_�_ �_o o2oDoVohozo �o�o�o�o�o�o�o
 .@Rdv�� �������*��<�N�`�r�������� ?��я�����+� =�O���r%{������� ß՟�����"�_���02�SwU�]n��� ������ȯگ���� "�4�F�X�j�|����� ��Ŀֿ�����0� B�T�f�xϊϜϮ��� ��������,�>ߩ� b�t߆ߘߪ߼����� ���o�(�:�L�^�p� �����#�Q�[�� ��
��.�@�R�d�v� �������������� '9K]o�� ������# 5GYk}�������O�3�/ /1/C/U/g/y/�/�/ �/�/�/�/�/	??-?�;:�D?q?{6���d�j?@]	12345678�R�h!B!�U���B��V� �?�?OO)O;OMO_O qOwA��O�O�O�O�O �O__*_<_N_`_r_ �_�_�_�_�]�O�_ o o$o6oHoZolo~o�o �o�o�o�o�o�o�_ �_DVhz��� ����
��.�@� R�d�#��������Џ ����*�<�N�`� r���������y�ޟ� ��&�8�J�\�n��� ������ȯگ���� ϟ4�F�X�j�|����� ��Ŀֿ�����0� B�T�f�%��ϜϮ��� ��������,�>�P� b�t߆ߘߪ߼�{��� ����(�:�L�^�p� ����������� ����0.�@�%����l�~����Cz � B\�   ���2d4� ���d1
���  	�d22,�%X7IXp���Z������� %7I[m �������� !/3/E/W/i/{/�/�/ �/�/�/�/�/??/?@A?S?e?w?�?�:Z������<�4��`�$�SCR_GRP �1�� �� � ���� ��	 _�1��2 
BD[����� I�7GpDO2OkO������hBDE� DP��wC�GhK�A�RC Mate �120iC 67w890��M-�@�A 8��M2I�A�A��
123�45�D;F�2  ����>U�1{F�1 HC�1�AhAJ<ANY	?R�_�_�_�_�_~�\��H��0�T�7�2 o/O0oVoho7F/��Co�o?o��o���l0Q�o:DB�B���r2tAA���A  @��YuA@9�Wpj ?�wr�H��DzAF@ F�`�r��o� ����B�-�f�Q� ��}Yq�r������ďքB��y�*��N� 9�r�]�o�����̟�� �۟�&���CTOF�k�����h�����q�Yq>��̣�7G@hYpݯ����W \HC+�3���AnpC�HV��o~ec��W���� y���������pո��¿ P�(�%�7�I�v�b�SS���0EL_DEFAULT  m�_���u�?HOTSTR�͐����MIPOWER�FL  ����޷�WFDO�� ��� u�RVENT? 1���`��� L!DUM�_EIPL�(��j�!AF_INEx��Fߺ�!FTߒu�<ߙ�!o�� ������!RP?C_MAIN����q���1���VIS���ٻ �}�!TP&p�PUt�/�dl����!
PMON_POROXY��2�e�������+�f�a�!�RDM_SRV�b�/�gP���!R�T��0�h����!
���M,�,�i��E!RLSYNCF�l	84�!R3OS߸�4���!
CE��MTC�OM�2�k�)!=	�CONS*1��lu!�WA'SRC|�2�md�;!�USB�0��n�/!STM��'/.�o�Y/��}/ p�J/\/�/�/�/�/���ICE_KL ?�%� (%S?VCPRG1�/::"$52:???)03b?g?")04�?�?)05�?�?")06�?�?)07OO�)0
TJOE<9ROWK &4��O)1,?�O)1T? �O)1|?�O)1�?_)1 �?G_)1�?o_)1O�_ )1DO�_)1lO�_Q1�O oQ1�O7oQ1�O_oQ1 _�oQ15_�oQ1]_�o Q1�_�oQ1�_'Q1�_ OQ1�_wy1%o�/	2 )0?"0���1�/� �S�>�w�b������� я��������=�(� a�L�s���������ߟ ʟ��'�9�$�]�H� ��l�����ɯ��ۯ�� �#��G�2�k�V��� ����ſ���Կ����1��C�g�Rϋ��*_�DEV ���MC:��t�����GRP 2��՟�0bx 	� 
 ,����ߟ���7��[� B�Tߑ�xߵߜ����� �����3�E�,�i�P� �������z������� ��A�S�:�w�^��� ������������+ O��D�<�� ����'9  ]D��z��� ��/h5/G/./k/ R/�/v/�/�/�/�/�/ ???C?*?g?y?`? �?�?�?�?*/�?�?O -OOQO8OuO�OnO�O �O�O�O�O_�O)__ M___F_�_�?x_�_p_ �_�_oo�_7oo[o moTo�oxo�o�o�o�o �o�oE�_i{ b������� ��A�S�:�w�^��� ����я�����^+� �O�a�H���l����� ��ߟƟ����9� � ]�D�����z������ �����5�G�.�k� R�������ſ����� ���C�*�<�yϟ�d ���	gϰϛ���Ͽ������+�%�x+�Pߌ����i� �i�y߇�qߧߕ��� ������=�"�e���O� =�s�a������� ��3��'��K�9�o� ]������������� ��#G5k��� ��[�W��� C�j�3�� �����/]B/ �/u/c/�/�/�/�/ �/�/5/?Y/�/M?;? q?_?�?�?�?�/�?�? �?�?�?OIO7OmO[O �O�?�O�?�O�O�O�O �O_E_3_i_�O�_�O Y_�_�_�_�_�_�_o Ao�_ho�_1o�o�o�o �o�o�o�oIooo@o sa����� !�E�9��I�o� ]��������ޏ��� ���5�#�E�k�Y��� я������ן��� 1��A�g�����͟W� �����ӯ	���-�o� T�f��?�������� �Ͽ�G�,�k���_� M�o�qσϹϧ���� �C���7�%�[�I�k� m�ߵ�����ߥ�� ��3�!�W�E�g���� ���ߍ��������/� �S���z���C���?� ��������+m�R ���s���� �E*i�]K �o����/ A�5/#/Y/G/}/k/ �/��/�/�/�/�/�/ 1??U?C?y?�/�?�/ i?�?�?�?�?�?-OO QO�?xO�?AO�O�O�O �O�O�O�O)_kOP_�O _�_q_�_�_�_�_�_ 1_W_(og_o[oIoo mo�o�o�o	o�o-o�o !�o1WE{i� �o������ -�S�A�w�����g� я�������)�O� ��v���?�����͟�� �ߟ�W�<�N��'� �o�����ɯ���/� �S�ݯG�5�W�Y�k� ����ſ��+���� �C�1�S�U�gϝ�߿ ��ύ������	�?� -�Oߥ��Ϝ���u��� ��������;�}�b� ��+��'������� ���U�:�y��m�[� �����������-� Q���E3iW�{ ���)� A/eS���� y�u�//=/+/ a/��/�Q/�/�/�/ �/�/??9?{/`?�/ )?�?�?�?�?�?�?�? OS?8Ow?OkOYO�O }O�O�O�OO?O_OO �OC_1_g_U_�_y_�_ �O�__�_	o�_o?o -ocoQo�o�_�o�_wo �o�o�o;)_ �o��oO���� ���7�y^��'� �������ُǏ��?� $�6����W���{� ����՟���;�ş/� �?�A�S���w���� ԯ������+��;� =�O���ǯ���u�߿ Ϳ��'��7ύ��� ��ÿ]Ϸϥ������� ��#�e�J߉��}�� �߳ߡ�������=�"� a���U�C�y�g��� �������9���-�� Q�?�u�c��������� �����)M; q����a�]� �%I�p� 9������� !/cH/�/{/i/�/ �/�/�/�/�/;/ ?_/ �/S?A?w?e?�?�?�? ?'?�?7?�?+OOOO =OsOaO�O�?�O�?�O �O�O_'__K_9_o_ �O�_�O__�_�_�_�_ �_#ooGo�_no�_7o �o�o�o�o�o�o�o aoF�oyg�� ���'���� �?�u�c�������� �#�����'�)�;� q�_���׏������� ݟ��#�%�7�m��� ��ӟ]�ǯ���ٯ� ���u���l���E��� ��ÿ���տ�M�2� q���e���uϛωϿ� ����%�
�I���=�+� a�O�qߗ߅߻����� !߫���9�'�]�K� m���ߺ��߃����� ���5�#�Y������ I�k�E��������� 1s�X��!�y� ����	K0o �cQ�u��� �#/G�;/)/_/ M/�/q/�/�/�// �/??7?%?[?I?? �/�?�/o?�?k?�?O �?3O!OWO�?~O�?GO �O�O�O�O�O_�O/_ qOV_�O_�_w_�_�_ �_�_�_oI_.om_�_ aoOo�oso�o�o�oo �o�o�o�o']K �o��o��� ���#�Y�G�}�� ���m�׏ŏ���� ��U���|���E��� ��ӟ������]��� T���-���u�����ϯ ���5��Y��M�߯ ]���q�����˿�� 1���%��I�7�Y�� mϣ����	ϓ����� !��E�3�U�{߽Ϣ� ��k����������� A��h�z�1�S�-�� ��������[�@������$SERV_MAIL  �����e�OUTP�UTt���RoV 2�	�  ��� (�O���i�S�AVE��g�TOP�10 2�� d ��;M_q ������� %7I[m� ������/!/ 3/E/W/i/{/�/�/�/ �/�/�/�/??/?	��YP��f�FZN_CFG �	�'��.��o1?GRP 2�y7��� ,B   A��0.D;� B��0�  B4.�RB21��HELLr2�	���������7"O1K%RSR1O2ODO}OhO�O �O�O�O�O�O�O_
_�C_._g_R_�_�_�^_�  ��%�_��_�_�R�\a. ��_b`ރ��R2�. do�_�6HK ;1��; o�o �o�o�o�o�o�o
3 .@R{v�������<OMM ���?2��2FTOV_ENBt�����HOW_REG_�UIR�g�IMIO/FWDL��!��5�A��*SYST�EM*. V8.3�0340 ł11�/9/2020 �A ���X��SNPX_ASG�_T   0 �$ADDRES�S  ��ZE��VAR_NAM�	�%$MULT�IPLY��P�ARAM�� � $TIME��v�$�_ID�	$NUM�D�T��CIMP[�FRI�FD�VERSIOyN��G�TATU ��$DISK�NF�OD�MODBUS�_ADR[�����P�ORC�۫�S�SR�� x =��NGLE��g��$DUMMY7��SGL�TASK   &�����T������STMyTT0�PSEGT2�BWD�h��E���SVCNT_G�P�� 8 $�PC�ER_V� �  	$FB:�Pm�SPC��m�� S�DX�R[��� �$DAT�A00�u���1���2��3��4��5���6��7��8��9���A��B��C��D��2���F�� y���U1Ω1۩1�1��U1�1�1�1)�U16�1C�1P�1]��1j�1w�ҀI���2�Ω2۩2�2��2��2�2�2)�2�6�2C�2P�2]�2�j�2w�3��3��3�Ω3۩3�3��3��3�3�3)�3�6�3C�3P�3]�3�j�3w�4��4��4�Ω4۩4�4��4��4�4�4)�4�6�4C�4P�4]�4�j�4w�5��5��5�Ω5۩5�5��5��5�5�5)�5�6�5C�5P�5]�5�j�5w�6��6��6�Ω6۩6�6��6��6�6�6)�6�6�6C�6P�6]�6�j�6w�7��7��7�Ω7۩7�7��7��7�7�7)�7�6�7C�7P�7]�7�j�7w�Q ��PR�M_UPDӑ � $4q� �
����ӑؐ$�TORQUE_C�MD   u�M}Oa_SPEEjQ_CURREo��nAXI �mS^�CART���_Ut��^/YS�LO� � ������������y_�{�VALU�COP��$�#(F��ID_L��K%HI�F*IN�$FI�LE_A�v$�$�M�t��SAR0 � h^� E_B�LCK���"���(D_CPU�)��)���F#y/�$���_=�R� 	 � P�WҐOT��)1LA#�SR� .3?184RUN_FLGQ58-4U184WITX5v1-4v185H2�D4�084�zg�TBC2���
 � $�O�X0IGu �0_F�TM1D��42D�T�DCX0AZ��2M0���6�1�7TH��C�DxGR.0A��ERVE�3?D�3?D�3O��0_AC@ X -$jA�LEN�3wD�3j@E�L_RATI��M$�W_�F#1jAc$2�GMO�!>��C>��ERTIA�o!0�Iaj@�KDE�E���LACEM�CC4�CmV�@MA��F87UW7QTCV>\_QWTRQ^\UuZ��`�Ct��USt�J_��q�M�TF�J2'���E)�QUvA2�P>��s�a�C@JKfV�K�1'a�1'a`A`J�0<d+cJJ3cJJ;cAAL+ca`3ca`�[f4\e5C�PN1��\�`Q[;P�L�@_��E�.�0CF�{ `^GROU1 (����y�N�0CC��`?REQUIR*B���EBUZ�fA�V$T�@2#qg@v�1�4 \�EN�ABL	�$AP�PRpCL�
$�OPEN`xCLO�SEozSE�y�E
\�1.� �u M�0p<PPB�t_MGr!�pC��� �x��9P�w�BRK�yNOLD|�vh�RTMO_�3H���uJ"��Pcd P3cP;cPcP�c�P6P��S�b� ��c�5� �r�B�1���1��PATH��ӁɃӁ�H�σ0�(p�W�SCaATr�ar�qINiB�UC�@��)�C��U%M2�Y�@+@�P9��O!EAT��0T�`@T�P�AYLOA�J2=L7R_AN�1���L*0���������uR_F2LSHR9DؑLO��(�ٗF��>F�ACRL_�!&���"���4bH$ ��$H�rG�FLEX�cs�0J�6 PMr�?�?>OPO�"d�>iE :vO�F P٧�O5aP�O�O�LF1�>�R��O�O �O�O_!_��E+_=_ O_a_s_�_�_�_�_Y� vĽW�Sdf����_�_H o�jT2'W�X� `�eŴ��e'� �*o <oNo``deme[ee�oКo�o�i�bJ�d ���0�o�o� 8A1Tk�q�PELٰ�1�=�xJ(p#pJE� �CTR"�f�TN�R9�wHAND_�VB�c�0 ��� $��F2�v	D�#SW���a�v� $$M���yv �q���q�����>���AR ���vQ!5��}A(�| �zA�{A�@��{� �zD�{D�P2�G@0��ST�w��4�y��N�DYW0^p �v!�H���k@ϗ�ϗ�ꑎ�g������P X�a�j�s�|��������ӵ5 ��Ť�����qASYM$��^�p������_�0�.�A�+��-��K�]�o�����J���K�����˙x�_�VI��	(�s V_UNIC.$P�בJeG"uG"�K$� X$|&
��P�K�,�>�$�%�T�\�\�a�0H+0Rr���!v�&VrDI�sO4��� �c `�O�I2AO�F�I1l�WW3�o��0�`ܰ�  o � ��ME���@r2�"YT0P�T���ڀ�1�`�d u���8�1�9T��a� $DUMM�Y1`A$PS_fi�RF+���$�6�XpFLA�`YP���B�3$GLB_T��5*E�0Vq�`8��j�v1 Xs�w֤�ST±#pSB}R��M21_VrT$SV_ER��1O� pC�CCLD@pBeAڰOL2� GL ;EW� 4�`�1W$YQ�ZQ�W�CH`ԑ��As02��"��@U�E ��N��@�$GIz�}$�A �@�C�@�� L�`V�}�$F�EVNEA�R��Np�F]Y��T�ANCp���JOG��A� ��$JOINT
Ѻ`�E�MSET�  "WECU۱�S�'U|��� g��U��?�#pLOC�K_FO���0B�GLVm�GLhT?EST_XMcp�Q'EMP�Pr+bBB��P$U���B2�2#p�CQab���PQarACE�`Sr`_ $KAR�M3TPDRA�@�d�Q�VEC��f�PIU�QaVaHE�PTO�OL2��cV1�REN�`IS3���b6s�Nf�ACH�P(p�a1O��3�429�2�`�ISr  @$R�AIL_BOXEz
��@ROBO"d�?��AHOWWA�RO�Aq�0qROLM�2gu��
txr��/p�Z���O_F��!� �D�a� �_ +�R�`Oˢ!�r*���Q�p�FOU�R"�XBMeYC���P/$PIP#fN���b�/r�ax�Qa�p��CORDED�P��q� ���OY0 # D )@OBu�G��P�d�S��3(@S��I�S;YSS�ADRH�� Κ0TCH�S� ,�0EN2�A�Q_�T������PVW�VAu1% � ��`�B5PREV�_RT�$ED�IT�VSHWRB��\F$����A	 �D�0��;���$HEAD�� U����KE�A�0CPwSPDl�JMPp��L5àR��44&�[�t���I,`SH�CƎ�NE�`I��TICK2�<M}����{HNRA' @]�8����t�_GP�&v΀�STY��qLO�DA�"����m�( �t 
 �Gƅ%$��T=\@S>�!�$=!2��1EF0FP�SQU�`%�B�!TERC�0Q�P��TS��)  Ph@�׹���g��a�`1O�0�3t�IZDQE�1PRE��1!�̯��pPU�1�_DYObR��XS�PK6�AXIP��sVaUR�ڳI�Hp�~����_�`��ET��P( bl�O�FP�A�4 ss�`��BSR��*lѠ��A����� ���#��1��A� R�c�R�s�RŃ�d�~� ��dŢ������ː́C��|����S}C,@ + h�@cDS��a�0SPC0&~�ATq��2������2ADDRESz�cB�SHIF�^H`_2CHH�z��IK@���TV�I�72,��h���� 
�+j
!P��>���- 	\����O����<�C��򢵲���B�<��TXSCRE�EU�.	0k�TICNA�CP��T�Q8����� / T���@ ����Ag@��^���^����RROL wP���f���h5�PUE��0# �� ��@S�A���RSM�T�UNEaX��6F�� S_�C�f�6V�i���6��Cx�RB��� 2/��UE�1=2�B��!�WGMT� Li!m�zw@O�WBBL_p9W�0��2 �O�5O�ALE���GpTO�3RIG�H&BRD�D��C�KGR�0NTEX���OJWIDTH@s1�u��1A�a%��I_�0H�� 3 8�!wP_T��ҭ�0R�@�Rsw�2$�R� O�ѭ�4���G�G U2 �R brqL�UM�u���ERV�
��@� PaP�У5z{0�GEUR&ciF���Q)]�LPM��E��C�)jS�xP�x�`w5u6u7u8Z���3�9�P��6�a�QS���4�USR�D6 <���0UR��R�FOC�aPPRI�αmp�!L TRI}P+qm�UN$0
547	Pt�$0��Yqp��Hb���� 8�\  �G \�T�p�1��ѣ"OS�1�&R ���#�a�9�O�C �N�"�$�IaUU��:�/�/�U��#OSFF!`��;[�3-On0 ٰW5�4�:�@GUNw�>�0B_SUB�2p@N��SRT� �<���vQ�p �ORp�5RAU��4T�9���19_���= |����OWN� T$S#RC���r�D!`CE�MPFI*�*ё�ESP-������e*�B�&�bE���>� `10WO8�T��COP:1$��� _^@�b�A�q�EWA�C?a�A�@�C8�A�b�PVCCH��? �qC36MFB1��R4�Y`��@x %rT���AXdP^��spC�p^RUDRIV���C_V�uT̐fpD�?MY_UBY�ZT V�񕠧�B��X�a��RP_Sp�+��RL�7�BM$��DEY��EX����E�MU��X7d[�UASP�po��G���PACINΑ}�RGMAadwbF3wb3wb���ARE����a�r�6Twb�pA R�@G"�PP�a6UR� �p�B d�_���2	l�BN�RECcSWo`�_Apa�8c�OD!��A��1s�E��UB�� �q5VHK
G�C��Iz���.p��zsEA���w�@� �1u5UMRCV��D� �FOS�M� C��	�rX3�c�rREF���v�v�q p7�� p �z��z��{;��vp_@@�zq��{���S�/g�Sᡏ�ѫ97S��E �$�=Џߠ) �UӠOU���b�ZS @�e2�2�$��R� �FΐB��2Ѻ�Kq��SUL�C�@C�O:�� D)`�NT�CZ��BY��e�!e�$�L�S���S���̚�!�JTǤFGt +��ǱT� ��oCACH+�LO�����*`����@ܣC�_LIMI��FR�%�Tj�'���$HO�� 6B�COMMpSB�O0 ]�Ԉ�I�؄h@VP�b��_'SZ3n���6����12���[`��&�����AaMP�FAIj&�Gvt��AD���BMREׄ9�_SIZ�PH�`��FASYNBUF�FVRTDk�w�I�a�OL��D_@3��W:3P�ETUc�yQNp[�ECCU�h�VEM�`��۲&�V�IRC���VTP��pO��J�s�A�w�_DELA�cP��Q�KS��G�p9pCKWLAS�3	ő_�$F�ƀHp"�S;��yN��PLEXEE�I��B/��4sFLK I `]�^A��M����dws3S/�^@�bJ# �ʱ��#�#RSn ORD@!���P> 3 ނ)�K���T\"���WwCb2V��g%L`�Qۑ6D�4��\*bUR4sp_R'�d���,a]��ծc �_od&�{g��`Br*�T�'�SCO��*�C� ad�"_f�"0� �">�"K�"Y�J_\_�nZ��� E\ AMܐP�0 PSM�f%Mp"%HADJ�T�/e��Bڒ� N8p"q׬!LIN]3q�/�XVRh$O\����T_OVR� �/ZABC�5P�bw�t$��
4QZIPg%}Qp"DBGLV�C�L�R ���MPCF�5R  r ���$���QLNK�2
8��-`|�S �|q��^��CMCMi`C�C�C�ACtP_�  �$J:4D ��@QJ�V�4p$0�tO�UXW� ��UXE>a��E��[���	��{�Z��T �����r�YK�D"0 �U�"��^IGHcq�?( �K���V � vG��$B$��@1e�BX�҉�&GRV%�F� ���OVC�5�A�7�w@�`��
VBI����D�TRAC�Ey V�1SPH�ER�P W ,� �3I[�$SI�M�A�!2Re!O� ��e!V&��qe!�8m/!��%���/Kp�b/t#_UN�@_+�p&LCд�% ��%V M��AL�IAS ?e����%1�! ( he�!:?L?^?p?�? �66?�?�?�?�?�?	O O-O?OQO�?uO�O�O �O�OhO�O�O__)_ �OM___q_�_._�_�_ �_�_�_�_o%o7oIo [ooo�o�o�o�oro �o�o!3�oWi {�8����� ��/�A�S�e���� ������я|����� +�֏<�a�s�����B� ��͟ߟ����'�9� K�]�o��������ɯ ۯ�����#�5��Y� k�}�����L�ſ׿� ��ϸ�1�C�U�g�y� $ϝϯ�����~���	� �-�?���c�u߇ߙ� ��V����������� ;�M�_�q��.��� �������%�7�I� ��m��������`��� ����!��EWi {&������ /AS�w� ���j��// +/�O/a/s/�/0/�/ �/�/�/�/�/?'?9?�K?]?3�$SMO�N_DEFPRO ����1� *SYSTEM*p:�RECALL ?�}�9 ( �}�:copy vi�rt:\outp�ut\untit�led1.pc �md: over� =>19175�8336:165�386d?O#O2K}�6�2frs:or�derfil.d�at�4tmpba�ck\�072.8�.9.225:7864 �?�O�O3O�-�2mdb:*.*[OmMtO__)_<F1xFD:\�OPP�OA �O�_�_�_@B2FUaN_`_�Cy_
oo.o AA�?�?�?�?�o�o�o� }
xyzra?te 11 Qoco uo*=E�g�[4092 �o�o����=Etpdi/sc 0P as���(�;Gtpc?onn 0 �� ��������o�aQ�c��u���*�=O}968�􏅟�����P� a�s���(�;�M� ݟ�������ɏ[��m���"�5�G�sB9756�����������P� a�s���(� ;�M�ܿ�2ϑϣ�6o�Ho�ol�88022�784:951580���#�6OHOZO R��ώߠ�3��O`�X� t���)�<_�_�_]� �߉����_Q�c�`� y�
��.�A�S����� ������������u� *=�����s�� �����^��& ���c������r=�F�rC132�P@dv//+/>�ƿ ����/�/�/<�N�@\/n/�/?#?6�7F��X�N/�P�/�?�?��. ��a?�u?OO*O�Ź3F?X8emp�L8�7`��?�O�O�O��+FF*.dZOlLsO_ _(_;�M��C�O�O�_ �_�_��R^a_s_oo (o�/M��_�_2o�o�o 6�HOZ?R^}o �o ���ooI�o�������$SNPX_A{SG������q�� P �0 '%R[1]@1.1��y?���%�(�� L�/�A���e������� ܏��я����H�+� l�O�a�������؟�� ��ߟ�2��<�h�K� ��o���¯��̯��ۯ ����R�5�\���k� �������ſ���� <��1�r�U�|Ϩϋ� �ϯ�������8�� \�?�Qߒ�uߜ��߫� ������"��,�X�;� |�_�q�������� ����B�%�L�x�[� ������������� ,!bEl�{ ������( L/A�e��� ���/�/H/+/ l/O/a/�/�/�/�/�/ �/�/�/2??<?h?K? �?o?�?�?�?�?�?�? O�?ORO5O\O�OkO �O�O�O�O�O�O_�O <__1_r_U_|_�_�_ �_�_�_o�_o8oo \o?oQo�ouo�o�o�d��tPARAM ��u�q ��	��jP;tAp��h#t��pOFT�_KB_CFG � s�u�sOPI�N_SIM  �{vu��p�p�RVQSTP_DSB^~r��x�`�SR ay �� & SOCgKET�"��v�TOP_ON_ERR  -�Kx?�_PTN �fr��A;�RIN�G_PRMI� ��`VCNT_GP� 2au&q�(px 	�̏p���ޏ���wVD��RP 1�i'p�y� R�d�v���������П �����*�<�N�`� ����������̯ޯ� ��&�M�J�\�n��� ������ȿڿ��� "�4�F�X�j�|ώϠ� ������������0� B�T�f�xߟߜ߮��� ��������,�>�e� b�t��������� ���+�(�:�L�^�p� ��������������  $6HZl~� ������  2DV}z��� ����
//C/@/ R/d/v/�/�/�/�/�/ �/	???*?<?N?`? r?�?�?�?�?�?�?�?�OO&O0�PRG_�COUN�At�8r�NuRBENB��ME�MwCAt�O_UPD� 1�{T  
;Or�O�O�O__ (_:_c_^_p_�_�_�_ �_�_�_�_ oo;o6o HoZo�o~o�o�o�o�o �o�o 2[V hz������ �
�3�.�@�R�{�v� ����Ï��Џ��� �*�S�N�`�r����� �����ޟ��+�&� 8�J�s�n��������� ȯگ����"�K�F� X�j���������ۿֿ ���#��0�B�k�f��x�DL_INFO {1�E�@��	 ����������>���@���j�������
� Aj������}�)L��S5�!և�Ad��o߁�� DlzD��Dh B���*��hx���*��ߤ�O@YSDOEBUG\@�@���d�I��SP_PA�SS\EB?��L_OG ���C����ؘ�  ���A��UD1:�\���_MPC �E���AH��� �Am�SAV ��m�4�L���S�SVd�TEM_TIME 1	�]�@ 0������)�[�L��$T1?SVGUNS�@]E�'�E�r�ASK_OPTION\@�E�A�A��_DI���xO��BC2_GRP 2
�I=���~��@�  C��CK��CFG ����� l�]`]`ߕ���� ���7"[F X�|����� �/3//W/B/{/f/ �/�/�/�/���,�/ �/"?4?�/?j?U?�? y?�?���?���0�? O �?$OOHO6OlOZO|O ~O�O�O�O�O�O_�O 2_ _B_h_V_�_z_�_ �_�_�_�_�_�_.oh � BoToro�o�oo�o �o�o�o�o&8 \J�n���� ���"��F�4�j� X�z�����ď���֏ �����0�f�T��� @o����ҟ���t�� �*�P�>�t�����f� �����ί���� (�^�L���p�����ʿ ��ڿ ��$��H�6� l�Z�|�~ϐ��ϴ��� ����2�D�V���z� hߊ߰ߞ��������� �
�@�.�d�R�t�v� �����������*� �:�`�N���r����� ����������&J  �bt���4� ���4FX& |j������ �//B/0/f/T/�/ x/�/�/�/�/�/?�/ ,??<?>?P?�?t?�? `�?�?�?OO�?:O (OJOpO^O�O�O�O�O �O�O _�O$__4_6_ H_~_l_�_�_�_�_�_ �_�_ ooDo2ohoVo �ozo�o�o�o�o�o
 �?"4Rdv�o� �������� <�*�`�N���r����� ��ޏ̏���&��J� 8�Z���n�����ȟ�� �ڟ�����F�4�j�  ������į֯T�����
�0��T�>�r���$TBCSG_G�RP 2>��  �r�� 
 ?�   ������ӿ������@-��Q�c�v�}����d0 ���?~r�	 HC�`��r���b�C�  B�����Ȣ�>�f�f�źƞ��������϶�\��H �h�BYLcφ�B$дh߀j߈ߎ߲߰����ތ��@�@��AƷ�f�y� D�V��������	�^�?333��2�	V3.00���	m2ia�	*T�L�q�c�"����r����� ���l���   ���B������u�J�2}���5���C�FG >���� ��
�D8��Go�o� �
G������ �5 YDV�z ������/1/ /U/@/y/d/�/�/�/ �/�/�/�/????Q? ����\?n?�?*?�?�? �?�?�?O�?1OOUO gOyO�OFO�O�O�O�O �O	_r�^�._:�>_@_ R_�_v_�_�_�_�_�_ �_o*ooNo<oro`o �o�o�o�o�o�o�o 8&\Jl�� ��������� 6�X�F�|�j�����ď ��ԏ����܏.�0� B�x�f�������ҟ�� �����*�,�>�t� b����������ί� ��:�(�^�L���p� ������ܿʿ ��$� �H�6�X�~�(��Ϩ� ��d����������D� 2�h�Vߌߞ߰��߀� ����
����@�R�d� �t��������� �����*�`�N��� r������������� &J8n\~� �����"�� :L
�|�� �����0/B/T/ /d/�/x/�/�/�/�/ �/?�/,??P?>?`? �?t?�?�?�?�?�?�? OOOLO:OpO^O�O �O�O�O�O�O�O_ _ 6_$_Z_H_j_l_~_�_ .�_�_�_�_ oo0o VoDozoho�o�o�o�o �o�o�o
@.P v��Tf��� ���<�*�L�r�`� ��������ޏ̏��� �8�&�\�J���n��� ����ڟȟ���"�� F�X�op���o>�į ���֯����B�0� f�x���H�Z������ ҿ��,�>���b�P� r�tφϼϪ������ ��(��8�^�L߂�p� �ߔ��߸�������$� �H�6�l�Z��~�� �����d����&��� ��D�V���z������� ����
.��R@ bdv����� �*N<^` r������/ /$/J/8/n/\/�/�/ �/�/�/�/�/?�/4? "?X?F?|?�?8��?�? �?t?�?�?OO.O0O BOxOfO�O�O�O�O�O��O�O__>_(^  9dPhS hV|_�hR�$TBJOP_GRP 20U��  �?�hV	�R�S��\�8P���p��Q�U � � � � y��RhS @dP��R	 �C� >ff  C�W�Q�4b��<f9o >��ff\a<a=�ZwC�`���b�&`H&`.g�o�g�nѴW4e\e`b�o �?a�d=�7LC��noBȂo#&`�p`9u�o�c�33\u�X2h�P<��C�\vc@333@�33|b}`�BL��wHqDa�l����u�Jh�p<X���B$�d��?_���C*p���C���Z`y�x��k<G ��q`?]`�C4.�ϏR�d��da�G����{<gș��]p@&b`yap�c�z{4ep�V� ���������ʟ��� (�� �N��Z����@������ޯ��d�hV�0�4e	V3.�00�Sm2ia�T*Z��TcQh�s�� E�'E��i�FV#F�"wqF>��F�Z� Fv�RF��~MF���F����F��=F����F�ъF���3F���F��{G
G�dG�G�#
��D���E'
EMK�E���E�ɑ�E�ۘE���E���F���F��F���F(��F5���FB��FO���F\��Fi���Fv��F��v�F�u�<#�
/<t���@Ť�Ar_X�j�M�hTn��@�U�S��SESTP�ARSA�\X�P�SH�R��ABLE 1%�[��hS�ȃ�Q �0cɞ����ȨgWoQ��	��
�������hQ����8��C���RDI�ϬQ��� �2�D�Vվ�O����������*���S�ߪS ������ �!�3�E�W�i�{��� ������������ /A�]�����̂	k� }���M�_�q߃ߕ������hNUM  �0U�Q�P�pP B�C���_CFGG P�a@�P�IMEBF_TT�����S���VER�AÔ��R 1=�[ 8e�hR�cP! 3P�   � //$/6/H/Z/l/ ~/�/�/�/�/�/�/�/ ? ?2?{?V?h?�?�? �?�?�?�?�>��?O�:0OBOTO.OxO�O dO�O�O�O�O�O�O_ ,__P_b_�8�_�_ �_~_�_�_�_�_����_K�@���M�I_CHAN� �� mcDBGLV�逡���p`ET�HERAD ?*���`�n��?o��o�o��p`ROUT6�!p
!"t@~|SNMASK�h|��a255.~u�F�|��F���OOLOFS_DI���GT �iORQC?TRL p	��	n��T�B�T�f� x���������ҏ��� ��,�>�P�b�r��𕟄�����PE_D�ETAI�h�zPG�L_CONFIG� Qa���/cell/$C�ID$/grp1���3�E�W�i�{�1� 	����ʯܯ� ��� $�6�H�Z�l�~���� ��ƿؿ�������2� D�V�h�zό�ϰ��� ������
ߙ�.�@�R� d�v߈��)߾���������}��N�`� r��������������)�;�M�_� �߃�����������l� %7I[m�� ������z !3EWi��� ������/// A/S/e/w//�/�/�/ �/�/�/�/?+?=?O? a?s?�??�?�?�?�? �?O�?'O9OKO]OoO �OO�O�O�O�O�O�O�_��User View !��}}1234567890B_T_f_x_��_�_�T-`��_��(Y25Y�Ooo*o<o No`o�_�_/R3�_�o �o�o�o�ogo)�^4�obt������^5Q�(�:�@L�^�p�����^6� ʏ܏� ��$���E��^7��~�������Ɵ؟7����^8m�2�D��V�h�z���럭��� �lCamera3Z)����(�:�L�*�E�v��� ��@_��ƿؿ�����  ̦�Y�^�p� �ϔϦϸ�_����� � K�$�6�H�Z�l�~ߥ��̦�i������� � �$���H�Z�l�ߐ� ���������ߣ�Py ��6�H�Z�l�~���7� ������#��� 2 DV���*����� ������"4F �j|����k ͥ��Y/ /2/D/V/ h/�/�/�/��/�/ �/
??.?���l��/ z?�?�?�?�?�?{/�? 
OOg?@OROdOvO�O �OA?�� �1O�O�O
_ _._@_�?d_v_�_�O �_�_�_�_�_o�O�G9�_GoYoko}o�o�o H_�o�o�o�_�o1�CUgy�	Υ0 �o�������o 2�D�V��oz������� ԏ{�Ӡիx�-� ?�Q�c�u���.����� ϟ����)�;�M� �ΥA�䟙�����ϯ �󯚟�)�;���_� q���������`��u�� P���)�;�M�_�� �ϕϧ��������� �%�̿޵���q߃� �ߧ߹���r����� ^�7�I�[�m���8� ޵�(�������%� 7���[�m������� ����������޵��� I[m��J�� ��6!3EW<i  	� �����//(/x:/L/^+   n v�/�/�/�/�/�/ ? ?$?6?H?Z?l?~?�? �?�?�?�?�?�?O O 2ODOVOhOzO�O�O�O �O�O�O�O
__._@_ R_d_v_�_�_�_�_�_�b,  
 (  ��( 	  �_oo:o(o^oLo�o po�o�o�o�o�o �ot$�Z~* ̸ i{� ���� ��X5�G�Y�� }�������ŏ׏��� ��f�C�U�g�y��� �����ӟ�,�	�� -�?�Q�c��������� �������)�;� ��_�q���ʯ����˿ ݿ��H�%�7�Iϐ� m�ϑϣϵ���� � ���!�h�E�W�i�{� �ߟ���������.�� �/�A�S�e�߉�� ������������+� r��a�s�������� ������J�'9K ��o����� ��X5GYk }������0 //1/C/U/g/��/ �/�/��/�/�/	?? -?t/Q?c?u?�/�?�?��?�?�?�?:?p@ AB"O4OFOCG� `��)frh:�\tpgl\ro�bots\m20�ia\arc_m�ate_1�@c.xmlO�O�O�O�O��O__(_:_L_XX��X_}_�_�_�_�_�_ �_�_oo1oCoZ_To yo�o�o�o�o�o�o�o 	-?VoPu� �������� )�;�RL�q������� ��ˏݏ���%�7� N�H�m��������ǟ ٟ����!�3�J�D� i�{�������ïկ� ����/�F�@�e�w� ��������ѿ������+�=�_H�1 �Oj@88�?�=�|�=�xϚϜ� ���������0��<� f�P�rߜ߆ߨ��߼�����&��$TPG�L_OUTPUT� "H1H1 `�H�]�o�� ������������� #�5�G�Y�k�}����������������H�`����2345678901 2DVh z�>2���� ��9K]o�}����� ���1/C/U/g/y/ �/#/�/�/�/�/�/	? �/???Q?c?u?�?? 1?�?�?�?�?OO�? %OMO_OqO�O�O-O�O �O�O�O__�O�OI_ [_m__�_�_;_�_�_ �_�_o!o�_/oWoio {o�o�o7oIo�o�o�o /�o=ew� ��E�����+�� �}[�a�s���������̍@b�����h� ( 	  7�%�[�I��m��� ������ǟ���!�� E�3�i�W�y�����ï ���կ�����/�e�S����^�w� ��ѽ�����)�;� ��d�v�ϚϬϊ� ����L���ߺ�(�N� ,�>߄ߖ� ߺ���n� �����&�8��D�n� �^��������V� �"���F�X�6�|��� ��z�����x����� 0B��fx�� ���N`,� Pb@���� p�/�/:/�� p/�/$/�/�/�/�/�/ X/�/$?�/4?Z?8?J? �?�??�?�?z?�?O �?2ODO�?POzOOjO �O�O�O�O�ObO_._ �OR_d_B_�_�__�_ �_�_�_oo�_<oNo�Tb�$TPOFF_LIM ���p�����qibNw_SVm`  ӄ�jP_MON �#���d�p��p2ӅiaSTRT?CHK $��f�^��bVTCOM�PAT�hq�fVW�VAR %�m\Ax�d �o Y��p�bia_DEFPROG 3v�b%SOCKE�p��m_DISP�LAYt`�n�rIN�ST_MSK  ��| �zINU�SER�tLCK���{QUICKM�ENA��tSCRE�`���rtpsc�t�{���b���_��STziR�ACE_CFG �&�iAtx`	�bt
?�܈HNL 2'�i}� �H{ nr4�F�X�j�|���𠟲�ĚޅITEM� 2( � �%�$1234567�890��  =�<�7�I�Q�  !W�_�kp���bs �ů)����_���� ��^���y�ݯ����5� %�7�I�c�m�翑�=� c�u�ٿ�����!ϛ� E����)ߍ�5߱��� ��Yߧ������A��� e�w�@��[���� �ߧ��k���O��s� �E�W���c������ }�'�����o�/�� ����;S����# �GY"}=�a s����1� U/'/����� �_/	/�/�/�/Q/? u/�/�/?�/i?�?�? ?�?)?;?M?�?O�? COUO�?aO�?�?�OO �O7O�O	_mO_�O�O l_�O�_�O�_�_�_3_ �_W_i_{_�_�_Koqo �o�_�ooo/o�o�o eo%7�oC�o�o� �o���O�s(�N�ڄS�)�S���  ϒS�q �����y
 ���ݏď���UD1�:\���e�R_�GRP 1*��� 	 @�p Y�k�U���y�����ӟ�������͑�2�x�V�A�?�  q� ��m�����ǯ���ٯ �����E�3�i�W���`{��������	!�����c�SCB 2+o� \�Y�k� }Ϗϡϳ�������Y��V_CONFIG ,o�󁧏�M����OUTPUT �-o�>��� Yߝ߯���������	� �-�?�Q�c�u�;ъ� �����������	�� -�?�Q�c�u������ ��������); M_q������ ��%7I[ m������ �/!/3/E/W/i/{/ ��/�/�/�/�/�/? ?/?A?S?e?w?�/�? �?�?�?�?�?OO+O =OOOaOsO�O�?�O�O �O�O�O__'_9_K_ ]_o_�_�O�_�_�_�_ �_�_o#o5oGoYoko }o�_�o�o�o�o�o�o 1CUgy� '�9Ո������ #�5�G�Y�k�}����� �oŏ׏�����1� C�U�g�y��������� ӟ���	��-�?�Q� c�u���������ϯ� ���)�;�M�_�q� ��������˿ݿ�� �%�7�I�[�m�ϑ� �ϴ����������!� 3�E�W�i�{ߍߟ߱� ����������/�A� S�e�w������� ������+�=�O�a� s��������������� '9K]o� �������� #5GYk}��|��x���� ���/�3/E/W/ i/{/�/�/�/�/�/�/ �/?�/?A?S?e?w? �?�?�?�?�?�?�?O O*?=OOOaOsO�O�O �O�O�O�O�O__&O 9_K_]_o_�_�_�_�_ �_�_�_�_o"_5oGo Yoko}o�o�o�o�o�o �o�o0oCUg y������� 	��,?�Q�c�u��� ������Ϗ���� (�;�M�_�q������� ��˟ݟ���%�6� I�[�m��������ǯ ٯ����!�2�E�W� i�{�������ÿտ������,��$TX�_SCREEN �1.����}ipnl�/`�gen.htm,�ϑϣϵ���$ �Panel �setup��}������0�B�T�f� ���ϝ߯��������� n���?�Q�c�u�� ���"��������� )�������q������� ����B���f�%7 I[m������� ���t��EW i{���:���////A/�/�U�ALRM_MSG� ?L��Y�  Z//��/�/�/�/�/�/ ??$?B?H?y?l?�?��?�?u%SEV  ��-�6s"EC�FG 0L��V�  /�@� � A#A   B�/�
 �?6�L�VO hOzO�O�O�O�O�O�O��O
_W�1GRP �21	K 0/�	� @Ob_u I_B�BL_NOTE �2	JT�G�l6�Q�8�@~uRDEFPRO =%�+ (%�?�_ 8��_o�_'ooKo6o ooZo�o�o�o�o�o�o�k\INUSER � �]P_�oI_M�ENHIST 1�3	I  ( ��P��(/SO�FTPART/G�ENLINK?c�urrent=m�enupage,153,17������)q�~381,23�/�A�S�2�'��~71������ӏ��q+y��ue�dit�rSOCKET��7�I�[��x���2���ȟڟ��r|p��148,2�>�P�b�t���o���� ��ϯ�󯂯�)�;� M�_�q�<x�Rlq��� ��Ϳ߿���'�9� K�]�oρ�ϥϷ��� �����ώϠ�5�G�Y� k�}ߏ�߳������� ����1�C�U�g�y� ���,���������	� ���?�Q�c�u����� ����������) ,�M_q���6 ���%7� [m���D� ��/!/3/�W/i/ {/�/�/�/�/R/�/�/ ??/?A?�/e?w?�? �?�?�?�����?OO +O=OOOR?sO�O�O�O �O�O\O�O__'_9_ K_]_�O�_�_�_�_�_ �_j_�_o#o5oGoYo �_}o�o�o�o�o�o�o xo1CUg�o �������?�? �-�?�Q�c�u�x�� ����Ϗ�󏂏��)� ;�M�_�q�������� ˟ݟ����%�7�I� [�m��� ���ǯٯ ������3�E�W�i� {������ÿտ��������$UI_�PANEDATA 15���A��  	��}  frh/�cgtp/wid�edev.stm��zόϞϰ���)  rih��ϧ�R� � �$�6�H�Z���lߐ� wߴߛ���������� 2�D�+�h�O������� � � �� � �����#�5�G�Y��� }��ϡ����������� b�1U<y� r�����	� -?&c���C� ��������P !/��E/W/i/{/�/�/ /�/�/�/�/�/?/? ?S?:?w?^?�?�?�? �?�?�?Oz�=OOO aOsO�O�O�?�O./�O �O__'_9_K_�Oo_ V_�_z_�_�_�_�_�_ o#o
oGo.oko}odo �oO&O�o�o�o 1�oUg�O��� ���L	��-�?� &�c�J����������� ��ڏ���;��o�o ~��������˟ݟ0� �t%�7�I�[�m�� 柣�����ٯ����� ��3��W�>�{���t� ����տ�Z�l��/� A�S�e�w�ʿ����� ��������+ߒ�O� 6�s�Zߗߩߐ��ߴ� �����'��K�]�D� ����Ϸ��������� �d�5�G���k�}��� ������,����� C*gy`�� ��������}�,ew����)S�W��/"/ 4/F/X/j/��/u/�/ �/�/�/�/?�/0?B? )?f?M?�?�?�?�?Q������$UI_P�OSTYPE  ���� �	 �?#O�2QU�ICKMEN  �KO&O�0RE�STORE 16���  '��?X��O�C�OX�m�O�O__'_ 9_�O]_o_�_�_�_H_ �_�_�_�_o�Oo0o Bo�_}o�o�o�o�oho �o�o1C�og y���Zo��� R�-�?�Q�c���� ������Ϗr���� )�;����Z�l�ޏ�� ��˟ݟ����%�7� I�[�m��������ǯ ٯ�����
�|�E�W� i�{���0���ÿտ� ��Ϯ�/�A�S�e�w��1GSCREA@?�FMu1sc��@u2��3��4���5��6��7��8<���2USER����2��T����ks���U4�5�6�7��8��0NDO_CFG 7K<;��0PDATE ���������4B��_INFO� 18����RA0%}���Q�������� '�
�K�]�@��d�� ����������*L���OFFSET ;FM�Ë@ �b� t��������������� N�UL^�� �����&VO(�
L*�UFRA_ME  �d����RTOL_AB�RTp�ӈENB���GRP 1<��IRACz  A������	//�-/?&I/[/�@@U��iѠMSK  ���ӢNm%��%��/�_EV�N��$c�
6U�2�=I9hi��UEV�!td�:\event_�user\�/T0C�7Y?)�F�<L1S�PR1W7spot�weld�=!CA6�?�?�?�@�$!�/ h?&O[OGl�OJO8O �O�OnO�O�O�O_�O �O�Oe__�_4_F_|_ �_�_�_�_�_�_=o,o aooo�oBo�o�oxo��o�o'�o�j)6W�RK 2>@�88"�� y�� ��
��.�@��d� v�Q�������Џ⏽� ���<�N�)�_���~���$VCCMUҳ?\ݨ�MR�2�E8;<�"�	�j���~XC5G6 *����h֜ �5�i�A@�7 p? ȗ� ;[�e�Ȇ���ů�����^�9%A���ٯ*�� B���E��I�ѯ j�����]�����ֿ�� �����0χ��f�Q��cϜ�O����ϥ�ISIONTMOU?� ��ů�FU���U�(�� FR:\��\�u�A�?  ��� MC*�LOG�7�   UD1�*�EX[�E!' B@ ���Ҁo�r���o������d ��  =	 �1- n6  G-����Ҭ6,��<��1�=���:����n�P�TRAI�N����1�E!�Adt��͓G8; (�� :��S����������� -��1�?�Q�c�u���Й���T���_��REⲐH�����LEX�E��I8;�1-e���VMPHASE'  ���A����RTD_FILT�ER 2J8; ��R����� ��1C#�� t��������//��SHIFT6�"1K8=<���/p/3��O/u/�/�/ �/�/�/�/?�/?)? b?9?K?�?o?�?�?�?�	LIVE/S�NAP�3vsf�liv4�?�>�� SETU�0BmenuOO�?}O��OfB/%L����	|H{O�O��?�J� ��@-�AdB8
�����K�M�QR��S����	'-_�ME�0�ļ�/!M�OM �zWqW�AITDINEN�D����TOK C 噰\���_S�_�YTIM����
lG�_,m�_Ok�_/j��_/jo�XRELE�K_g���Q��֗Q_�ACT�0^h(q�X_N3� N��)r%�Ox_��rRDIS�0~�n�$XVR�B�O �$ZABCv͒1P�� ,��r��2g7ZIP�CQ����/�A�S��z�MPCF_G 1	R�J�0��w��a��MP�sS���<������8��?Vv����>�t�
t��? �?Z����p�C�d�>���DlzD�Dh���?��>������*�=E������4�X>C�����"�4�;B�T�f����Ο�����A�2�B��*��?hx��*�*�<�>ȿߐn�h�z�����ȫ�pt��T|��w�_YLINDqU|��  �e� ,(  *)�:���&�c�J���n� ���Ͽ �#��s�(��!�^� ���ϔϦ����e�K�  ���$��y�Z�l��{���2V�+q � ���������������٧�D��ז^�A����SPHERE 2W	�̾Ϛ�ߓ� �����<�O�*�<��� `������}������ ��I�[�8��\C�U�������pZZ�f ��f