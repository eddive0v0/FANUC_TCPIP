��   ��A��*SYST�EM*��V8.3�0340 11�/9/2020 A 	  ����PASSNA�ME_T   �0 $+ �$'WORD � ? LEVEL � $TI- OUTT  &F/�� $SE�TUPJPROG�RAMJINST�ALLJY  $CURR_OަUSER�NU�M�STPS_L�OG_P N��$��T�N�  �6 COUNT_D�OWN�$EN�B_PCMPWD� � DV�I�N!$C� C{RE�PARM:z� T:DIAG:�)�LVCHK|!FULLM0�YXT�CNTyD�MENU��AUTO,�FG�_DSP�RLS��U�&ENC�/  C�RYPTE  }1�$$CL(   ���;!��� D 0 V� IO�� :&  ���L!IRTU�A� :/�$DCSo_COD@���?%�  W�'_WS  v*�!x ��&�A91�"w!{� 
 $B! ���-�/? ?6?D?Z? h?~?�?�?�?�?�?�?��?OO2O���#SUP� �+4OFO�#F�fOxO�O�� � �L�A���O �� �� V�[_t&��j���D�ON_��W
_��d ��V�U�YWALUGH� 1w) d �)�_�_�_o o)o;oMo_oqo�o�o �o�'�_�o�o�o /ASew��� �o�����+�=� O�a�s��������� ߏ���'�9�K�]� o���������Ə۟� ���#�5�G�Y�k�}� ������¯���� �1�C�U�g�y����� ����Я���	��-� ?�Q�c�uχϙϫϽ� ̿������)�;�M� _�q߃ߕߧ߹����� ����%�7�I�[�m� ������������ �!�3�E�W�i�{��� ������������ /ASew��� ���%