��  I��A��*SYST�EM*��V8.3�0340 11�/9/2020 A   ����SBR_T �  | 	$S�VMTR_ID � $ROBO�T9$GRP�_NUM<AXIaSQ6K 6NFF�3 _PARAM�F	$�  �,$MD SPD�_LIT  &2�*� � ��  �$$CLA�SS  ���������� V�ERSION��  ��~�IRTUAL���'  1 �� T���A�RC Mate �120iC���  �aiS12�/4000 80�A��
H1 D�SP1-S1��	P01.05W,  	� v���  ��# :�����������{  ���r9 � �9����� HH��  �����
/ms��� D4�~Z %%������ ����� 1�2M���?�X���B=�d������&���<
= z ����� J����������; �� � ���T����N�.����Y	� � � !� ��� :�?8���'by�c/�/�/�/L?��?;?!�R?d?v?�?��2/�1��>��x����r�߼2*->�0�����o��G>�?�?��<RN`r2|2�j� ���  J � 	������,������A �'/�/��A#�"p<� 2�"t��=���	��7�_��
��D<)�J � ����� EV$���?p$��z(>�]�q"��P�(�/ �/���/�_�_�_�_ ?��_D?oo1oCo�0��"��@����
�P,$bb�3dH�@~������:3�#uFo�o�T�?N�@8Nw3�|3<ONI
[K&�����wB
�=� �D���S�J8HB �,P����.��+ ]^'H�H�&�����1�/���>���� � �23
��K>vB� ��
P�@�X"��op# ��Z{ 2|%j��`R� ��l�&W�BVR� d^Sco A�jS:rY:q�K�]�o� ���_�����ҏ���`��,�>���ɬo�Nb@/6
!A4�k4|b�o����P��ϓ�p�`�M������{��9�9� ���"�@D@o�r� ���X"��  ��'��sBC�U����/ 	����,V$y����  �� �z�s;@2��q"��� �D�_%���p(����'jT�rYT����� '�9���]���������@��ɿۿ���Z��d�.N��R��x�5|�b��Ԛ�������X� � �/X"��  �!-�?��������*�p$q�P�r�1�ϾzR��Q ��&� į֯诱�������B� �f�/�A�S�e�w������N@�r6|6d�v�О=����Ҩ��k ��2�X"��Q��������-�8����t ��!�����qTa
��#�&�|ߎߠ�i{� ��������/ASew�����xTa���Ng�	�LA ���/ /2/D/V/ h/z/�/�/�/�/�/�/@�/
??.?@?P<�P? t?�?�?�?�?�?�?�? OO(O0C��FO� ���O�O�O�O�O_ _*_<_N_`_r_�_�_ �_�_�_�_�_o^?&o 8oJo\ono�o�o�o�o �o�o6OhOZO#~O�O Xj|����� ����0�B�T�f� x�������
o����� ��,�>�P�b�t��� ���o����*<N� (�:�L�^�p������� ��ʯܯ� ��$�6� H�Z�l�ȏ������ƿ ؿ���� �2�D�V� ҟğn��������� ��
��.�@�R�d�v� �ߚ߬߾�������� �*N�`�r��� ����������^ϐ� ��K��ϸπ������� ��������"4F Xj|����� 2��0BTf x������� R�d�v�>/P/b/t/�/ �/�/�/�/�/�/?? (?:?L?^?p?�?�?� �?�?�?�? OO$O6O HOZOlO~O���O/ "/4/�O_ _2_D_V_ h_z_�_�_�_�_�_�_ �_
oo.o@oRo�?vo �o�o�o�o�o�o�o *�O�O�Os�O�O �������&� 8�J�\�n��������� ȏڏ���Zo�4�F� X�j�|�������ğ֟ �D� �z��f� x���������ү��� ��,�>�P�b�t��� ����������� (�:�L�^�pςϔϦ� "����8�J�\�$�6� H�Z�l�~ߐߢߴ��� ������� �2�D�V� h�z�ֿ��������� ��
��.�@�R����� �ϛ���������� *<N`r�� �����& ��8\n���� ����/l�5/(/ �������/�/�/�/�/ �/�/??0?B?T?f? x?�?�?�?�?�?�?@ OO,O>OPObOtO�O �O�O�O�OJ/</�O`/ r/�/L_^_p_�_�_�_ �_�_�_�_ oo$o6o HoZolo~o�o�o�?�o �o�o�o 2DV hz�O_�O�_0_ �
��.�@�R�d�v� ��������Џ��� �*�<�N��o`����� ����̟ޟ���&� 8��]�P������ ȯگ����"�4�F� X�j�|�������Ŀֿ ����h�0�B�T�f� xϊϜϮ��������� r�d�߈�����t߆� �ߪ߼��������� (�:�L�^�p���� ����&��� ��$�6� H�Z�l�~�������0� "���F�X� 2DV hz������ �
.@Rdv �������/ /*/</N/`/���/x/ ���/�/??&? 8?J?\?n?�?�?�?�? �?�?�?�?O"O4O� XOjO|O�O�O�O�O�O �O�O__�/�/6_�/ �/�/�_�_�_�_�_�_ oo,o>oPoboto�o �o�o�o�o�o�oNO (:L^p��� ��&_X_J_�n_�_ H�Z�l�~�������Ə ؏���� �2�D�V� h�z������o��ԟ� ��
��.�@�R�d�v� ��������,�>�� �*�<�N�`�r����� ����̿޿���&� 8�J�\ϸ��ϒϤ϶� ���������"�4�F� ¯��^�د������� ������0�B�T�f� x������������ ��v�>�P�b�t��� ������������N߀� r�;�ߨ�p��� ���� $6 HZl~���� "���/ /2/D/V/ h/z/�/�/�/�/�/ BTf.?@?R?d?v? �?�?�?�?�?�?�?O O*O<ONO`OrO�O� �O�O�O�O�O__&_ 8_J_\_n_�/�/�_ ? ?$?�_�_o"o4oFo Xojo|o�o�o�o�o�o �o�o0B�Of x������� ��v_�_�_c��_�_ ������Ώ����� (�:�L�^�p������� ��ʟܟ�J �$�6� H�Z�l�~�������Ư د4����j�|���V� h�z�������¿Կ� ��
��.�@�R�d�v� �ϚϬ��������� �*�<�N�`�r߄ߖ� ����(�:�L��&� 8�J�\�n����� ���������"�4�F� X�j��ώ��������� ����0B���� �ߋ�������� ,>Pbt� ������// r�(/L/^/p/�/�/�/ �/�/�/�/ ?\%?? ���~?�?�?�?�? �?�?�?O O2ODOVO hOzO�O�O�O�O�O0/ �O
__._@_R_d_v_ �_�_�_�_:?,?�_P? b?t?<oNo`oro�o�o �o�o�o�o�o& 8J\n���O� �����"�4�F� X�j��_�_�_��o o �����0�B�T�f� x���������ҟ��� ��,�>��P�t��� ������ί���� (���M�@���̏ޏ�� ��ʿܿ� ��$�6� H�Z�l�~ϐϢϴ��� ������X� �2�D�V� h�zߌߞ߰������� b�T���x�����d�v� ������������ �*�<�N�`�r����� ���������& 8J\n���� � ��6�H�"4F Xj|����� ��//0/B/T/f/ ��x/�/�/�/�/�/�/ ??,?>?P?�u?h? ���?�?�?OO (O:OLO^OpO�O�O�O �O�O�O�O __$_�/ H_Z_l_~_�_�_�_�_ �_�_�_o�?|?&o�? �?�?�o�o�o�o�o�o �o
.@Rdv ������>_� �*�<�N�`�r����� ����oHo:o�^opo 8�J�\�n��������� ȟڟ����"�4�F� X�j�|������į֯ �����0�B�T�f� x�ԏ����
��.��� ��,�>�P�b�tφ� �Ϫϼ��������� (�:�Lߨ�p߂ߔߦ� �������� ��$�6� ����N�ȿڿ쿴��� ������� �2�D�V� h�z������������� ��
f�.@Rdv ������>�p� b�+���`r�� �����//&/ 8/J/\/n/�/�/�/�/ �/�/�/?"?4?F? X?j?|?�?�?��?�? 2DVO0OBOTOfO xO�O�O�O�O�O�O�O __,_>_P_b_t_�/ �_�_�_�_�_�_oo (o:oLo^o�?�?vo�? OO�o�o $6 HZl~���� ���� �2��_V� h�z�������ԏ� ��
�fo�o�oS��o�o ��������П���� �*�<�N�`�r����� ����̯ޯ:���&� 8�J�\�n��������� ȿ$���Z�l�~�F� X�j�|ώϠϲ����� ������0�B�T�f� xߊߜ����������� ��,�>�P�b�t�� ������*�<��� (�:�L�^�p������� �������� $6 HZ��~���� ��� 2���� ��{������� �
//./@/R/d/v/ �/�/�/�/�/�/�/? b?<?N?`?r?�?�? �?�?�?�?�?LOO ���nO�O�O�O�O �O�O�O�O_"_4_F_ X_j_|_�_�_�_�_ ? �_�_oo0oBoTofo xo�o�o�o*OO�o@O ROdO,>Pbt� �������� (�:�L�^�p����_�� ��ʏ܏� ��$�6� H�Z��o�o�o���o ؟���� �2�D�V� h�z�������¯ԯ� ��
��.���@�d�v� ��������п���� �t�=�0Ϫ���Ο�� �Ϻ���������&� 8�J�\�n߀ߒߤ߶� ������H��"�4�F� X�j�|�������� R�D���h�zό�T�f� x��������������� ,>Pbt� ������ (:L^p���� ��&�8� //$/6/ H/Z/l/~/�/�/�/�/ �/�/�/? ?2?D?V? �h?�?�?�?�?�?�? �?
OO.O@O�eOXO ����O�O�O�O_ _*_<_N_`_r_�_�_ �_�_�_�_�_oop? 8oJo\ono�o�o�o�o �o�o�o�ozOlO�O �O�O|����� ����0�B�T�f� x���������ҏ.o�� ��,�>�P�b�t��� ����8*�N` (�:�L�^�p������� ��ʯܯ� ��$�6� H�Z�l�~�ڏ����ƿ ؿ���� �2�D�V� h�ğ�π������� ��
��.�@�R�d�v� �ߚ߬߾�������� �*�<`�r��� �����������&� �ϔ�>������Ϥ��� ��������"4F Xj|����� ��V�0BTf x�����.�`� R�/v���P/b/t/�/ �/�/�/�/�/�/?? (?:?L?^?p?�?�?�? �?�?�? OO$O6O HOZOlO~O�O��O�O "/4/F/_ _2_D_V_ h_z_�_�_�_�_�_�_ �_
oo.o@oRodo�? �o�o�o�o�o�o�o *<N�O�Of�O �O_�����&� 8�J�\�n��������� ȏڏ����"�~oF� X�j�|�������ğ֟ ���V�zC��� x���������ү��� ��,�>�P�b�t��� ������ο*���� (�:�L�^�pςϔϦ� �������J�\�n�6� H�Z�l�~ߐߢߴ��� ������� �2�D�V� h�z��述������� ��
��.�@�R�d�v� ���ώ���,��� *<N`r�� �����& 8J��n���� ����/"/~��� ��k/�����/�/�/�/ �/�/??0?B?T?f? x?�?�?�?�?�?�?�? RO,O>OPObOtO�O �O�O�O�O�O</_�O r/�/�/^_p_�_�_�_ �_�_�_�_ oo$o6o HoZolo~o�o�o�oO �o�o�o 2DV hz��__�0_ B_T_�.�@�R�d�v� ��������Џ��� �*�<�N�`�r��o�� ����̟ޟ���&� 8�J������� � ȯگ����"�4�F� X�j�|�������Ŀֿ �����z�0�T�f� xϊϜϮ��������� �d�-� ߚ������� �ߪ߼��������� (�:�L�^�p���� ������8� ��$�6� H�Z�l�~��������� B�4���X�j�|�DV hz������ �
.@Rdv �������/ /*/</N/`/r/��  ���/(�/??&? 8?J?\?n?�?�?�?�? �?�?�?�?O"O4OFO �XO|O�O�O�O�O�O �O�O__0_�/U_H_ �/�/�/�_�_�_�_�_ oo,o>oPoboto�o �o�o�o�o�o�o`O (:L^p��� ����j_\_��_ �_�_l�~�������Ə ؏���� �2�D�V� h�z�������� ��
��.�@�R�d�v� �����(���>�P� �*�<�N�`�r����� ����̿޿���&� 8�J�\�n�ʟ�Ϥ϶� ���������"�4�F� Xߴ�}�p������� ������0�B�T�f� x������������ ��,���P�b�t��� ������������ �߄�.�ߺ��ߔ� ���� $6 HZl~���� ��F�/ /2/D/V/ h/z/�/�/�/�/P B?fx@?R?d?v? �?�?�?�?�?�?�?O O*O<ONO`OrO�O�O ��O�O�O�O__&_�8_J_\_n_�_�%�$SBR2 1 5��P T0 ��  @?7  �_�_�_o o2oDoVo hozo�o�o�o�o�o�Q �o�_ 2DVh z������� �o��o@�R�d�v��� ������Џ���� *��N�1�r������� ��̟ޟ���&�8� J�\�?���c�����ȯ گ����"�4�F�X� j�|���q�����ֿ� ����0�B�T�f�x� �ϜϮ��ϣ�~�_�� ���!�3�E�W�i�{� �ߟ߱����������� �(�:�L�^�p��� ��������� ���� �H�Z�l�~������� �������� 2D (�:�z����� ��
.@Rd vZ������ //*/</N/`/r/�/ �/�/��/�/�/?? &?8?J?\?n?�?�?�? �?�?�?�/�?O"O4O FOXOjO|O�O�O�O�O �O�O�O_�?0_B_T_ f_x_�_�_�_�_�_�_ �_oo,o>o"_boto �o�o�o�o�o�o�o (:L^pTo� ����� ��$� 6�H�Z�l�~������ Ə؏���� �2�D� V�h�z��������� ����
��.�@�R�d� v���������Я��� ؟�*�<�N�`�r��� ������̿޿��� &�
�4�\�nπϒϤ� �����������"�4� F�X�<�|ߎߠ߲��� ��������0�B�T� f�x��n߮������� ����,�>�P�b�t� �������������� (:L^p�� �������$ 6HZl~��� ����/ /D/ V/h/z/�/�/�/�/�/ �/�/
??.?@?R?6/ v?�?�?�?�?�?�?�? OO*O<ONO`OrOV? h?�O�O�O�O�O__ &_8_J_\_n_�_�_�_ �O�O�_�_�_o"o4o FoXojo|o�o�o�o�o �o�_�o0BT fx������ ���o,�>�P�b�t� ��������Ώ���� �(�:��^�p����� ����ʟܟ� ��$� 6�H�Z�l�P������� Ưد���� �2�D� V�h�z�������¿Կ ���
��.�@�R�d� vψϚϬϾ��ϴ��� ��*�<�N�`�r߄� �ߨߺ���������� &�8�J�\�n���� �����������"�� �X�j�|��������� ������0BT 8�J������� �,>Pbt �j�����/ /(/:/L/^/p/�/�/ �/�/��/�/ ??$? 6?H?Z?l?~?�?�?�? �?�?�?�/O O2ODO VOhOzO�O�O�O�O�O �O�O
__ O@_R_d_ v_�_�_�_�_�_�_�_ oo*o<oNo2_ro�o �o�o�o�o�o�o &8J\n�do� ������"�4� F�X�j�|�������� ֏�����0�B�T� f�x���������ҟ�� ȏ��,�>�P�b�t� ��������ί��� ���:�L�^�p����� ����ʿܿ� ��$� 6��D�l�~ϐϢϴ� ��������� �2�D� V�h�Lόߞ߰����� ����
��.�@�R�d� v���~߾������� ��*�<�N�`�r��� ������������ &8J\n��� �������"4 FXj|���� ���//0/T/ f/x/�/�/�/�/�/�/ �/??,?>?P?b?F/ �?�?�?�?�?�?�?O O(O:OLO^OpO�Of? x?�O�O�O�O __$_ 6_H_Z_l_~_�_�_�_ �O�O�_�_o o2oDo Vohozo�o�o�o�o�o �o�_�o.@Rd v������� ���o<�N�`�r��� ������̏ޏ���� &�8�J�.�n������� ��ȟڟ����"�4� F�X�j�|�`�����į ֯�����0�B�T� f�x���������ҿ� ����,�>�P�b�t� �ϘϪϼ�����Ŀ� �(�:�L�^�p߂ߔ� �߸������� ���� 6�H�Z�l�~���� ��������� �2�� (�h�z����������� ����
.@Rd H�Z������� *<N`r� �z����// &/8/J/\/n/�/�/�/ �/�/��/�/?"?4? F?X?j?|?�?�?�?�? �?�?�?�/O0OBOTO fOxO�O�O�O�O�O�O �O__,_OP_b_t_ �_�_�_�_�_�_�_o o(o:oLo^oB_�o�o �o�o�o�o�o $ 6HZl~�to� ����� �2�D� V�h�z�������� ���
��.�@�R�d� v���������П�Ə ؏�*�<�N�`�r��� ������̯ޯ��� ��
�J�\�n������� ��ȿڿ����"�4� F�*�T�|ώϠϲ��� ��������0�B�T� f�x�\Ϝ߮������� ����,�>�P�b�t� ������������ �(�:�L�^�p����� ���������� $ 6HZl~��� ������2D Vhz����� ��
//./@/$d/ v/�/�/�/�/�/�/�/ ??*?<?N?`?r?V/ �?�?�?�?�?�?OO &O8OJO\OnO�O�Ov? �?�O�O�O�O_"_4_ F_X_j_|_�_�_�_�_ �O�O�_oo0oBoTo foxo�o�o�o�o�o�o �o�_,>Pbt �������� �(�L�^�p����� ����ʏ܏� ��$� 6�H�Z�l�